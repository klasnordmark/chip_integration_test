VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_io
  CLASS BLOCK ;
  FOREIGN chip_io ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1758.200 32.990 1820.800 95.440 ;
    END
  END clock
  PIN clock_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.635 208.565 1756.915 210.965 ;
    END
  END clock_core
  PIN analog_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.705 4977.035 718.985 4979.435 ;
    END
  END analog_en[0]
  PIN analog_pol[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.265 4977.035 712.545 4979.435 ;
    END
  END analog_pol[0]
  PIN analog_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.085 4977.035 697.365 4979.435 ;
    END
  END analog_sel[0]
  PIN dm[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.485 4977.035 715.765 4979.435 ;
    END
  END dm[0]
  PIN dm[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.685 4977.035 724.965 4979.435 ;
    END
  END dm[1]
  PIN dm[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.865 4977.035 694.145 4979.435 ;
    END
  END dm[2]
  PIN enh[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.065 4977.035 703.345 4979.435 ;
    END
  END enh[0]
  PIN hldh_n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.845 4977.035 700.125 4979.435 ;
    END
  END hldh_n[0]
  PIN holdover[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.645 4977.035 690.925 4979.435 ;
    END
  END holdover[0]
  PIN ib_mode_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.465 4977.035 675.745 4979.435 ;
    END
  END ib_mode_sel[0]
  PIN inp_dis[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.505 4977.035 709.785 4979.435 ;
    END
  END inp_dis[0]
  PIN io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 679.200 5092.560 741.800 5155.010 ;
    END
  END io[0]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.085 4977.035 743.365 4979.435 ;
    END
  END io_in[0]
  PIN io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.885 4977.035 688.165 4979.435 ;
    END
  END io_out[0]
  PIN oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.245 4977.035 672.525 4979.435 ;
    END
  END oeb[0]
  PIN slow_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.885 4977.035 734.165 4979.435 ;
    END
  END slow_sel[0]
  PIN vtrip_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.685 4977.035 678.965 4979.435 ;
    END
  END vtrip_sel[0]
  PIN analog_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 782.705 210.965 782.985 ;
    END
  END analog_en[10]
  PIN analog_pol[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 776.265 210.965 776.545 ;
    END
  END analog_pol[10]
  PIN analog_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 761.085 210.965 761.365 ;
    END
  END analog_sel[10]
  PIN dm[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 779.485 210.965 779.765 ;
    END
  END dm[30]
  PIN dm[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 788.685 210.965 788.965 ;
    END
  END dm[31]
  PIN dm[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 757.865 210.965 758.145 ;
    END
  END dm[32]
  PIN enh[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 767.065 210.965 767.345 ;
    END
  END enh[10]
  PIN hldh_n[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 763.845 210.965 764.125 ;
    END
  END hldh_n[10]
  PIN holdover[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 754.645 210.965 754.925 ;
    END
  END holdover[10]
  PIN ib_mode_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 739.465 210.965 739.745 ;
    END
  END ib_mode_sel[10]
  PIN inp_dis[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 773.505 210.965 773.785 ;
    END
  END inp_dis[10]
  PIN io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 743.200 95.440 805.800 ;
    END
  END io[10]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 807.085 210.965 807.365 ;
    END
  END io_in[10]
  PIN io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 751.885 210.965 752.165 ;
    END
  END io_out[10]
  PIN oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 736.245 210.965 736.525 ;
    END
  END oeb[10]
  PIN slow_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 797.885 210.965 798.165 ;
    END
  END slow_sel[10]
  PIN vtrip_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 742.685 210.965 742.965 ;
    END
  END vtrip_sel[10]
  PIN analog_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1391.705 210.965 1391.985 ;
    END
  END analog_en[11]
  PIN analog_pol[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1385.265 210.965 1385.545 ;
    END
  END analog_pol[11]
  PIN analog_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1370.085 210.965 1370.365 ;
    END
  END analog_sel[11]
  PIN dm[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1388.485 210.965 1388.765 ;
    END
  END dm[33]
  PIN dm[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1397.685 210.965 1397.965 ;
    END
  END dm[34]
  PIN dm[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1366.865 210.965 1367.145 ;
    END
  END dm[35]
  PIN enh[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1376.065 210.965 1376.345 ;
    END
  END enh[11]
  PIN hldh_n[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1372.845 210.965 1373.125 ;
    END
  END hldh_n[11]
  PIN holdover[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1363.645 210.965 1363.925 ;
    END
  END holdover[11]
  PIN ib_mode_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1348.465 210.965 1348.745 ;
    END
  END ib_mode_sel[11]
  PIN inp_dis[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1382.505 210.965 1382.785 ;
    END
  END inp_dis[11]
  PIN io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1352.200 95.440 1414.800 ;
    END
  END io[11]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1416.085 210.965 1416.365 ;
    END
  END io_in[11]
  PIN io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1360.885 210.965 1361.165 ;
    END
  END io_out[11]
  PIN oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1345.245 210.965 1345.525 ;
    END
  END oeb[11]
  PIN slow_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1406.885 210.965 1407.165 ;
    END
  END slow_sel[11]
  PIN vtrip_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1351.685 210.965 1351.965 ;
    END
  END vtrip_sel[11]
  PIN analog_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1999.705 210.965 1999.985 ;
    END
  END analog_en[12]
  PIN analog_pol[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1993.265 210.965 1993.545 ;
    END
  END analog_pol[12]
  PIN analog_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1978.085 210.965 1978.365 ;
    END
  END analog_sel[12]
  PIN dm[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1996.485 210.965 1996.765 ;
    END
  END dm[36]
  PIN dm[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2005.685 210.965 2005.965 ;
    END
  END dm[37]
  PIN dm[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1974.865 210.965 1975.145 ;
    END
  END dm[38]
  PIN enh[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1984.065 210.965 1984.345 ;
    END
  END enh[12]
  PIN hldh_n[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1980.845 210.965 1981.125 ;
    END
  END hldh_n[12]
  PIN holdover[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1971.645 210.965 1971.925 ;
    END
  END holdover[12]
  PIN ib_mode_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1956.465 210.965 1956.745 ;
    END
  END ib_mode_sel[12]
  PIN inp_dis[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1990.505 210.965 1990.785 ;
    END
  END inp_dis[12]
  PIN io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1960.200 95.440 2022.800 ;
    END
  END io[12]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2024.085 210.965 2024.365 ;
    END
  END io_in[12]
  PIN io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1968.885 210.965 1969.165 ;
    END
  END io_out[12]
  PIN oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1953.245 210.965 1953.525 ;
    END
  END oeb[12]
  PIN slow_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2014.885 210.965 2015.165 ;
    END
  END slow_sel[12]
  PIN vtrip_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1959.685 210.965 1959.965 ;
    END
  END vtrip_sel[12]
  PIN analog_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2608.705 210.965 2608.985 ;
    END
  END analog_en[13]
  PIN analog_pol[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2602.265 210.965 2602.545 ;
    END
  END analog_pol[13]
  PIN analog_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2587.085 210.965 2587.365 ;
    END
  END analog_sel[13]
  PIN dm[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2605.485 210.965 2605.765 ;
    END
  END dm[39]
  PIN dm[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2614.685 210.965 2614.965 ;
    END
  END dm[40]
  PIN dm[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2583.865 210.965 2584.145 ;
    END
  END dm[41]
  PIN enh[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2593.065 210.965 2593.345 ;
    END
  END enh[13]
  PIN hldh_n[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2589.845 210.965 2590.125 ;
    END
  END hldh_n[13]
  PIN holdover[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2580.645 210.965 2580.925 ;
    END
  END holdover[13]
  PIN ib_mode_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2565.465 210.965 2565.745 ;
    END
  END ib_mode_sel[13]
  PIN inp_dis[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2599.505 210.965 2599.785 ;
    END
  END inp_dis[13]
  PIN io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2569.200 95.440 2631.800 ;
    END
  END io[13]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2633.085 210.965 2633.365 ;
    END
  END io_in[13]
  PIN io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2577.885 210.965 2578.165 ;
    END
  END io_out[13]
  PIN oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2562.245 210.965 2562.525 ;
    END
  END oeb[13]
  PIN slow_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2623.885 210.965 2624.165 ;
    END
  END slow_sel[13]
  PIN vtrip_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2568.685 210.965 2568.965 ;
    END
  END vtrip_sel[13]
  PIN analog_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3217.705 210.965 3217.985 ;
    END
  END analog_en[14]
  PIN analog_pol[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3211.265 210.965 3211.545 ;
    END
  END analog_pol[14]
  PIN analog_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3196.085 210.965 3196.365 ;
    END
  END analog_sel[14]
  PIN dm[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3214.485 210.965 3214.765 ;
    END
  END dm[42]
  PIN dm[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3223.685 210.965 3223.965 ;
    END
  END dm[43]
  PIN dm[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3192.865 210.965 3193.145 ;
    END
  END dm[44]
  PIN enh[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3202.065 210.965 3202.345 ;
    END
  END enh[14]
  PIN hldh_n[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3198.845 210.965 3199.125 ;
    END
  END hldh_n[14]
  PIN holdover[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3189.645 210.965 3189.925 ;
    END
  END holdover[14]
  PIN ib_mode_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3174.465 210.965 3174.745 ;
    END
  END ib_mode_sel[14]
  PIN inp_dis[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3208.505 210.965 3208.785 ;
    END
  END inp_dis[14]
  PIN io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3178.200 95.440 3240.800 ;
    END
  END io[14]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3242.085 210.965 3242.365 ;
    END
  END io_in[14]
  PIN io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3186.885 210.965 3187.165 ;
    END
  END io_out[14]
  PIN oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3171.245 210.965 3171.525 ;
    END
  END oeb[14]
  PIN slow_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3232.885 210.965 3233.165 ;
    END
  END slow_sel[14]
  PIN vtrip_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3177.685 210.965 3177.965 ;
    END
  END vtrip_sel[14]
  PIN analog_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3825.705 210.965 3825.985 ;
    END
  END analog_en[15]
  PIN analog_pol[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3819.265 210.965 3819.545 ;
    END
  END analog_pol[15]
  PIN analog_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3804.085 210.965 3804.365 ;
    END
  END analog_sel[15]
  PIN dm[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3822.485 210.965 3822.765 ;
    END
  END dm[45]
  PIN dm[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3831.685 210.965 3831.965 ;
    END
  END dm[46]
  PIN dm[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3800.865 210.965 3801.145 ;
    END
  END dm[47]
  PIN enh[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3810.065 210.965 3810.345 ;
    END
  END enh[15]
  PIN hldh_n[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3806.845 210.965 3807.125 ;
    END
  END hldh_n[15]
  PIN holdover[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3797.645 210.965 3797.925 ;
    END
  END holdover[15]
  PIN ib_mode_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3782.465 210.965 3782.745 ;
    END
  END ib_mode_sel[15]
  PIN inp_dis[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3816.505 210.965 3816.785 ;
    END
  END inp_dis[15]
  PIN io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3786.200 95.440 3848.800 ;
    END
  END io[15]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3850.085 210.965 3850.365 ;
    END
  END io_in[15]
  PIN io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3794.885 210.965 3795.165 ;
    END
  END io_out[15]
  PIN oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3779.245 210.965 3779.525 ;
    END
  END oeb[15]
  PIN slow_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3840.885 210.965 3841.165 ;
    END
  END slow_sel[15]
  PIN vtrip_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3785.685 210.965 3785.965 ;
    END
  END vtrip_sel[15]
  PIN analog_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.705 4977.035 1263.985 4979.435 ;
    END
  END analog_en[1]
  PIN analog_pol[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.265 4977.035 1257.545 4979.435 ;
    END
  END analog_pol[1]
  PIN analog_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.085 4977.035 1242.365 4979.435 ;
    END
  END analog_sel[1]
  PIN dm[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.485 4977.035 1260.765 4979.435 ;
    END
  END dm[3]
  PIN dm[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.685 4977.035 1269.965 4979.435 ;
    END
  END dm[4]
  PIN dm[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.865 4977.035 1239.145 4979.435 ;
    END
  END dm[5]
  PIN enh[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.065 4977.035 1248.345 4979.435 ;
    END
  END enh[1]
  PIN hldh_n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.845 4977.035 1245.125 4979.435 ;
    END
  END hldh_n[1]
  PIN holdover[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.645 4977.035 1235.925 4979.435 ;
    END
  END holdover[1]
  PIN ib_mode_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.465 4977.035 1220.745 4979.435 ;
    END
  END ib_mode_sel[1]
  PIN inp_dis[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.505 4977.035 1254.785 4979.435 ;
    END
  END inp_dis[1]
  PIN io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1224.200 5092.560 1286.800 5155.010 ;
    END
  END io[1]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.085 4977.035 1288.365 4979.435 ;
    END
  END io_in[1]
  PIN io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.885 4977.035 1233.165 4979.435 ;
    END
  END io_out[1]
  PIN oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.245 4977.035 1217.525 4979.435 ;
    END
  END oeb[1]
  PIN slow_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.885 4977.035 1279.165 4979.435 ;
    END
  END slow_sel[1]
  PIN vtrip_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.685 4977.035 1223.965 4979.435 ;
    END
  END vtrip_sel[1]
  PIN analog_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.705 4977.035 1808.985 4979.435 ;
    END
  END analog_en[2]
  PIN analog_pol[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.265 4977.035 1802.545 4979.435 ;
    END
  END analog_pol[2]
  PIN analog_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.085 4977.035 1787.365 4979.435 ;
    END
  END analog_sel[2]
  PIN dm[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.485 4977.035 1805.765 4979.435 ;
    END
  END dm[6]
  PIN dm[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1814.685 4977.035 1814.965 4979.435 ;
    END
  END dm[7]
  PIN dm[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.865 4977.035 1784.145 4979.435 ;
    END
  END dm[8]
  PIN enh[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.065 4977.035 1793.345 4979.435 ;
    END
  END enh[2]
  PIN hldh_n[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.845 4977.035 1790.125 4979.435 ;
    END
  END hldh_n[2]
  PIN holdover[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.645 4977.035 1780.925 4979.435 ;
    END
  END holdover[2]
  PIN ib_mode_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.465 4977.035 1765.745 4979.435 ;
    END
  END ib_mode_sel[2]
  PIN inp_dis[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.505 4977.035 1799.785 4979.435 ;
    END
  END inp_dis[2]
  PIN io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1769.200 5092.560 1831.800 5155.010 ;
    END
  END io[2]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1833.085 4977.035 1833.365 4979.435 ;
    END
  END io_in[2]
  PIN io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.885 4977.035 1778.165 4979.435 ;
    END
  END io_out[2]
  PIN oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.245 4977.035 1762.525 4979.435 ;
    END
  END oeb[2]
  PIN slow_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.885 4977.035 1824.165 4979.435 ;
    END
  END slow_sel[2]
  PIN vtrip_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.685 4977.035 1768.965 4979.435 ;
    END
  END vtrip_sel[2]
  PIN analog_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.705 4977.035 2353.985 4979.435 ;
    END
  END analog_en[3]
  PIN analog_pol[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2347.265 4977.035 2347.545 4979.435 ;
    END
  END analog_pol[3]
  PIN analog_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2332.085 4977.035 2332.365 4979.435 ;
    END
  END analog_sel[3]
  PIN dm[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2359.685 4977.035 2359.965 4979.435 ;
    END
  END dm[10]
  PIN dm[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.865 4977.035 2329.145 4979.435 ;
    END
  END dm[11]
  PIN dm[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.485 4977.035 2350.765 4979.435 ;
    END
  END dm[9]
  PIN enh[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2338.065 4977.035 2338.345 4979.435 ;
    END
  END enh[3]
  PIN hldh_n[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.845 4977.035 2335.125 4979.435 ;
    END
  END hldh_n[3]
  PIN holdover[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.645 4977.035 2325.925 4979.435 ;
    END
  END holdover[3]
  PIN ib_mode_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.465 4977.035 2310.745 4979.435 ;
    END
  END ib_mode_sel[3]
  PIN inp_dis[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.505 4977.035 2344.785 4979.435 ;
    END
  END inp_dis[3]
  PIN io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2314.200 5092.560 2376.800 5155.010 ;
    END
  END io[3]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.085 4977.035 2378.365 4979.435 ;
    END
  END io_in[3]
  PIN io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.885 4977.035 2323.165 4979.435 ;
    END
  END io_out[3]
  PIN oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.245 4977.035 2307.525 4979.435 ;
    END
  END oeb[3]
  PIN slow_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.885 4977.035 2369.165 4979.435 ;
    END
  END slow_sel[3]
  PIN vtrip_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.685 4977.035 2313.965 4979.435 ;
    END
  END vtrip_sel[3]
  PIN analog_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 757.015 3379.435 757.295 ;
    END
  END analog_en[4]
  PIN analog_pol[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 763.455 3379.435 763.735 ;
    END
  END analog_pol[4]
  PIN analog_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 778.635 3379.435 778.915 ;
    END
  END analog_sel[4]
  PIN dm[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 760.235 3379.435 760.515 ;
    END
  END dm[12]
  PIN dm[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 751.035 3379.435 751.315 ;
    END
  END dm[13]
  PIN dm[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 781.855 3379.435 782.135 ;
    END
  END dm[14]
  PIN enh[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 772.655 3379.435 772.935 ;
    END
  END enh[4]
  PIN hldh_n[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 775.875 3379.435 776.155 ;
    END
  END hldh_n[4]
  PIN holdover[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 785.075 3379.435 785.355 ;
    END
  END holdover[4]
  PIN ib_mode_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 800.255 3379.435 800.535 ;
    END
  END ib_mode_sel[4]
  PIN inp_dis[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 766.215 3379.435 766.495 ;
    END
  END inp_dis[4]
  PIN io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 734.200 3555.010 796.800 ;
    END
  END io[4]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 732.635 3379.435 732.915 ;
    END
  END io_in[4]
  PIN io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 787.835 3379.435 788.115 ;
    END
  END io_out[4]
  PIN oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 803.475 3379.435 803.755 ;
    END
  END oeb[4]
  PIN slow_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 741.835 3379.435 742.115 ;
    END
  END slow_sel[4]
  PIN vtrip_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 797.035 3379.435 797.315 ;
    END
  END vtrip_sel[4]
  PIN analog_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1366.015 3379.435 1366.295 ;
    END
  END analog_en[5]
  PIN analog_pol[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1372.455 3379.435 1372.735 ;
    END
  END analog_pol[5]
  PIN analog_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1387.635 3379.435 1387.915 ;
    END
  END analog_sel[5]
  PIN dm[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1369.235 3379.435 1369.515 ;
    END
  END dm[15]
  PIN dm[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1360.035 3379.435 1360.315 ;
    END
  END dm[16]
  PIN dm[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1390.855 3379.435 1391.135 ;
    END
  END dm[17]
  PIN enh[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1381.655 3379.435 1381.935 ;
    END
  END enh[5]
  PIN hldh_n[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1384.875 3379.435 1385.155 ;
    END
  END hldh_n[5]
  PIN holdover[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1394.075 3379.435 1394.355 ;
    END
  END holdover[5]
  PIN ib_mode_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1409.255 3379.435 1409.535 ;
    END
  END ib_mode_sel[5]
  PIN inp_dis[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1375.215 3379.435 1375.495 ;
    END
  END inp_dis[5]
  PIN io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1343.200 3555.010 1405.800 ;
    END
  END io[5]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1341.635 3379.435 1341.915 ;
    END
  END io_in[5]
  PIN io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1396.835 3379.435 1397.115 ;
    END
  END io_out[5]
  PIN oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1412.475 3379.435 1412.755 ;
    END
  END oeb[5]
  PIN slow_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1350.835 3379.435 1351.115 ;
    END
  END slow_sel[5]
  PIN vtrip_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1406.035 3379.435 1406.315 ;
    END
  END vtrip_sel[5]
  PIN analog_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1974.015 3379.435 1974.295 ;
    END
  END analog_en[6]
  PIN analog_pol[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1980.455 3379.435 1980.735 ;
    END
  END analog_pol[6]
  PIN analog_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1995.635 3379.435 1995.915 ;
    END
  END analog_sel[6]
  PIN dm[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1977.235 3379.435 1977.515 ;
    END
  END dm[18]
  PIN dm[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1968.035 3379.435 1968.315 ;
    END
  END dm[19]
  PIN dm[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1998.855 3379.435 1999.135 ;
    END
  END dm[20]
  PIN enh[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1989.655 3379.435 1989.935 ;
    END
  END enh[6]
  PIN hldh_n[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1992.875 3379.435 1993.155 ;
    END
  END hldh_n[6]
  PIN holdover[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2002.075 3379.435 2002.355 ;
    END
  END holdover[6]
  PIN ib_mode_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2017.255 3379.435 2017.535 ;
    END
  END ib_mode_sel[6]
  PIN inp_dis[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1983.215 3379.435 1983.495 ;
    END
  END inp_dis[6]
  PIN io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1951.200 3555.010 2013.800 ;
    END
  END io[6]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1949.635 3379.435 1949.915 ;
    END
  END io_in[6]
  PIN io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2004.835 3379.435 2005.115 ;
    END
  END io_out[6]
  PIN oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2020.475 3379.435 2020.755 ;
    END
  END oeb[6]
  PIN slow_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1958.835 3379.435 1959.115 ;
    END
  END slow_sel[6]
  PIN vtrip_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2014.035 3379.435 2014.315 ;
    END
  END vtrip_sel[6]
  PIN analog_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2583.015 3379.435 2583.295 ;
    END
  END analog_en[7]
  PIN analog_pol[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2589.455 3379.435 2589.735 ;
    END
  END analog_pol[7]
  PIN analog_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2604.635 3379.435 2604.915 ;
    END
  END analog_sel[7]
  PIN dm[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2586.235 3379.435 2586.515 ;
    END
  END dm[21]
  PIN dm[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2577.035 3379.435 2577.315 ;
    END
  END dm[22]
  PIN dm[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2607.855 3379.435 2608.135 ;
    END
  END dm[23]
  PIN enh[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2598.655 3379.435 2598.935 ;
    END
  END enh[7]
  PIN hldh_n[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2601.875 3379.435 2602.155 ;
    END
  END hldh_n[7]
  PIN holdover[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2611.075 3379.435 2611.355 ;
    END
  END holdover[7]
  PIN ib_mode_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2626.255 3379.435 2626.535 ;
    END
  END ib_mode_sel[7]
  PIN inp_dis[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2592.215 3379.435 2592.495 ;
    END
  END inp_dis[7]
  PIN io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2560.200 3555.010 2622.800 ;
    END
  END io[7]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2558.635 3379.435 2558.915 ;
    END
  END io_in[7]
  PIN io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2613.835 3379.435 2614.115 ;
    END
  END io_out[7]
  PIN oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2629.475 3379.435 2629.755 ;
    END
  END oeb[7]
  PIN slow_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2567.835 3379.435 2568.115 ;
    END
  END slow_sel[7]
  PIN vtrip_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2623.035 3379.435 2623.315 ;
    END
  END vtrip_sel[7]
  PIN analog_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3192.015 3379.435 3192.295 ;
    END
  END analog_en[8]
  PIN analog_pol[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3198.455 3379.435 3198.735 ;
    END
  END analog_pol[8]
  PIN analog_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3213.635 3379.435 3213.915 ;
    END
  END analog_sel[8]
  PIN dm[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3195.235 3379.435 3195.515 ;
    END
  END dm[24]
  PIN dm[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3186.035 3379.435 3186.315 ;
    END
  END dm[25]
  PIN dm[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3216.855 3379.435 3217.135 ;
    END
  END dm[26]
  PIN enh[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3207.655 3379.435 3207.935 ;
    END
  END enh[8]
  PIN hldh_n[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3210.875 3379.435 3211.155 ;
    END
  END hldh_n[8]
  PIN holdover[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3220.075 3379.435 3220.355 ;
    END
  END holdover[8]
  PIN ib_mode_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3235.255 3379.435 3235.535 ;
    END
  END ib_mode_sel[8]
  PIN inp_dis[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3201.215 3379.435 3201.495 ;
    END
  END inp_dis[8]
  PIN io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3169.200 3555.010 3231.800 ;
    END
  END io[8]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3167.635 3379.435 3167.915 ;
    END
  END io_in[8]
  PIN io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3222.835 3379.435 3223.115 ;
    END
  END io_out[8]
  PIN oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3238.475 3379.435 3238.755 ;
    END
  END oeb[8]
  PIN slow_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3176.835 3379.435 3177.115 ;
    END
  END slow_sel[8]
  PIN vtrip_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3232.035 3379.435 3232.315 ;
    END
  END vtrip_sel[8]
  PIN analog_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3800.015 3379.435 3800.295 ;
    END
  END analog_en[9]
  PIN analog_pol[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3806.455 3379.435 3806.735 ;
    END
  END analog_pol[9]
  PIN analog_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3821.635 3379.435 3821.915 ;
    END
  END analog_sel[9]
  PIN dm[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3803.235 3379.435 3803.515 ;
    END
  END dm[27]
  PIN dm[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3794.035 3379.435 3794.315 ;
    END
  END dm[28]
  PIN dm[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3824.855 3379.435 3825.135 ;
    END
  END dm[29]
  PIN enh[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3815.655 3379.435 3815.935 ;
    END
  END enh[9]
  PIN hldh_n[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3818.875 3379.435 3819.155 ;
    END
  END hldh_n[9]
  PIN holdover[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3828.075 3379.435 3828.355 ;
    END
  END holdover[9]
  PIN ib_mode_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3843.255 3379.435 3843.535 ;
    END
  END ib_mode_sel[9]
  PIN inp_dis[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3809.215 3379.435 3809.495 ;
    END
  END inp_dis[9]
  PIN io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3777.200 3555.010 3839.800 ;
    END
  END io[9]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3775.635 3379.435 3775.915 ;
    END
  END io_in[9]
  PIN io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3830.835 3379.435 3831.115 ;
    END
  END io_out[9]
  PIN oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3846.475 3379.435 3846.755 ;
    END
  END oeb[9]
  PIN slow_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3784.835 3379.435 3785.115 ;
    END
  END slow_sel[9]
  PIN vtrip_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3840.035 3379.435 3840.315 ;
    END
  END vtrip_sel[9]
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1226.430 4954.040 1226.750 4954.100 ;
        RECT 1352.470 4954.040 1352.790 4954.100 ;
        RECT 1572.810 4954.040 1573.130 4954.100 ;
        RECT 1226.430 4953.900 1352.790 4954.040 ;
        RECT 1226.430 4953.840 1226.750 4953.900 ;
        RECT 1352.470 4953.840 1352.790 4953.900 ;
        RECT 1545.760 4953.900 1573.130 4954.040 ;
        RECT 681.330 4953.700 681.650 4953.760 ;
        RECT 1448.610 4953.700 1448.930 4953.760 ;
        RECT 1545.760 4953.700 1545.900 4953.900 ;
        RECT 1572.810 4953.840 1573.130 4953.900 ;
        RECT 1573.270 4954.040 1573.590 4954.100 ;
        RECT 1573.270 4953.900 1642.040 4954.040 ;
        RECT 1573.270 4953.840 1573.590 4953.900 ;
        RECT 681.330 4953.560 1090.500 4953.700 ;
        RECT 681.330 4953.500 681.650 4953.560 ;
        RECT 1090.360 4953.360 1090.500 4953.560 ;
        RECT 1448.610 4953.560 1476.440 4953.700 ;
        RECT 1448.610 4953.500 1448.930 4953.560 ;
        RECT 1476.300 4953.360 1476.440 4953.560 ;
        RECT 1476.760 4953.560 1545.900 4953.700 ;
        RECT 1641.900 4953.700 1642.040 4953.900 ;
        RECT 1641.900 4953.560 1642.500 4953.700 ;
        RECT 1476.760 4953.360 1476.900 4953.560 ;
        RECT 1090.360 4953.220 1186.640 4953.360 ;
        RECT 1476.300 4953.220 1476.900 4953.360 ;
        RECT 1642.360 4953.360 1642.500 4953.560 ;
        RECT 1862.610 4953.360 1862.930 4953.420 ;
        RECT 2316.630 4953.360 2316.950 4953.420 ;
        RECT 2318.010 4953.360 2318.330 4953.420 ;
        RECT 1642.360 4953.220 1642.960 4953.360 ;
        RECT 1186.500 4953.020 1186.640 4953.220 ;
        RECT 1226.430 4953.020 1226.750 4953.080 ;
        RECT 1186.500 4952.880 1226.750 4953.020 ;
        RECT 1642.820 4953.020 1642.960 4953.220 ;
        RECT 1862.610 4953.220 2318.330 4953.360 ;
        RECT 1862.610 4953.160 1862.930 4953.220 ;
        RECT 2316.630 4953.160 2316.950 4953.220 ;
        RECT 2318.010 4953.160 2318.330 4953.220 ;
        RECT 1766.470 4953.020 1766.790 4953.080 ;
        RECT 1642.820 4952.880 1766.790 4953.020 ;
        RECT 1226.430 4952.820 1226.750 4952.880 ;
        RECT 1766.470 4952.820 1766.790 4952.880 ;
        RECT 1766.470 4951.660 1766.790 4951.720 ;
        RECT 1771.530 4951.660 1771.850 4951.720 ;
        RECT 1862.610 4951.660 1862.930 4951.720 ;
        RECT 1766.470 4951.520 1862.930 4951.660 ;
        RECT 1766.470 4951.460 1766.790 4951.520 ;
        RECT 1771.530 4951.460 1771.850 4951.520 ;
        RECT 1862.610 4951.460 1862.930 4951.520 ;
        RECT 2318.010 4950.440 2318.330 4950.700 ;
        RECT 2318.100 4950.300 2318.240 4950.440 ;
        RECT 3367.270 4950.300 3367.590 4950.360 ;
        RECT 2318.100 4950.160 3367.590 4950.300 ;
        RECT 3367.270 4950.100 3367.590 4950.160 ;
        RECT 3367.270 3839.520 3367.590 3839.580 ;
        RECT 3376.930 3839.520 3377.250 3839.580 ;
        RECT 3367.270 3839.380 3377.250 3839.520 ;
        RECT 3367.270 3839.320 3367.590 3839.380 ;
        RECT 3376.930 3839.320 3377.250 3839.380 ;
        RECT 208.910 3786.480 209.230 3786.540 ;
        RECT 212.590 3786.480 212.910 3786.540 ;
        RECT 208.910 3786.340 212.910 3786.480 ;
        RECT 208.910 3786.280 209.230 3786.340 ;
        RECT 212.590 3786.280 212.910 3786.340 ;
        RECT 3367.730 3726.640 3368.050 3726.700 ;
        RECT 3376.010 3726.640 3376.330 3726.700 ;
        RECT 3367.730 3726.500 3376.330 3726.640 ;
        RECT 3367.730 3726.440 3368.050 3726.500 ;
        RECT 3376.010 3726.440 3376.330 3726.500 ;
        RECT 213.050 3238.880 213.370 3239.140 ;
        RECT 213.140 3238.740 213.280 3238.880 ;
        RECT 213.140 3238.600 213.740 3238.740 ;
        RECT 212.130 3237.720 212.450 3237.780 ;
        RECT 213.600 3237.720 213.740 3238.600 ;
        RECT 212.130 3237.580 213.740 3237.720 ;
        RECT 212.130 3237.520 212.450 3237.580 ;
        RECT 3367.730 3231.600 3368.050 3231.660 ;
        RECT 3376.930 3231.600 3377.250 3231.660 ;
        RECT 3367.730 3231.460 3377.250 3231.600 ;
        RECT 3367.730 3231.400 3368.050 3231.460 ;
        RECT 3376.930 3231.400 3377.250 3231.460 ;
        RECT 212.130 3215.280 212.450 3215.340 ;
        RECT 213.510 3215.280 213.830 3215.340 ;
        RECT 212.130 3215.140 213.830 3215.280 ;
        RECT 212.130 3215.080 212.450 3215.140 ;
        RECT 213.510 3215.080 213.830 3215.140 ;
        RECT 208.910 3178.560 209.230 3178.620 ;
        RECT 211.210 3178.560 211.530 3178.620 ;
        RECT 213.510 3178.560 213.830 3178.620 ;
        RECT 208.910 3178.420 213.830 3178.560 ;
        RECT 208.910 3178.360 209.230 3178.420 ;
        RECT 211.210 3178.360 211.530 3178.420 ;
        RECT 213.510 3178.360 213.830 3178.420 ;
        RECT 210.750 3091.520 211.070 3091.580 ;
        RECT 211.670 3091.520 211.990 3091.580 ;
        RECT 210.750 3091.380 211.990 3091.520 ;
        RECT 210.750 3091.320 211.070 3091.380 ;
        RECT 211.670 3091.320 211.990 3091.380 ;
        RECT 210.750 3090.840 211.070 3090.900 ;
        RECT 211.670 3090.840 211.990 3090.900 ;
        RECT 210.750 3090.700 211.990 3090.840 ;
        RECT 210.750 3090.640 211.070 3090.700 ;
        RECT 211.670 3090.640 211.990 3090.700 ;
        RECT 210.750 2994.960 211.070 2995.020 ;
        RECT 212.130 2994.960 212.450 2995.020 ;
        RECT 210.750 2994.820 212.450 2994.960 ;
        RECT 210.750 2994.760 211.070 2994.820 ;
        RECT 212.130 2994.760 212.450 2994.820 ;
        RECT 212.130 2898.060 212.450 2898.120 ;
        RECT 213.050 2898.060 213.370 2898.120 ;
        RECT 212.130 2897.920 213.370 2898.060 ;
        RECT 212.130 2897.860 212.450 2897.920 ;
        RECT 213.050 2897.860 213.370 2897.920 ;
        RECT 212.130 2801.500 212.450 2801.560 ;
        RECT 213.510 2801.500 213.830 2801.560 ;
        RECT 212.130 2801.360 213.830 2801.500 ;
        RECT 212.130 2801.300 212.450 2801.360 ;
        RECT 213.510 2801.300 213.830 2801.360 ;
        RECT 213.510 2787.560 213.830 2787.620 ;
        RECT 213.970 2787.560 214.290 2787.620 ;
        RECT 213.510 2787.420 214.290 2787.560 ;
        RECT 213.510 2787.360 213.830 2787.420 ;
        RECT 213.970 2787.360 214.290 2787.420 ;
        RECT 3367.730 2617.900 3368.050 2617.960 ;
        RECT 3376.930 2617.900 3377.250 2617.960 ;
        RECT 3367.730 2617.760 3377.250 2617.900 ;
        RECT 3367.730 2617.700 3368.050 2617.760 ;
        RECT 3376.930 2617.700 3377.250 2617.760 ;
        RECT 208.910 2574.380 209.230 2574.440 ;
        RECT 211.670 2574.380 211.990 2574.440 ;
        RECT 213.510 2574.380 213.830 2574.440 ;
        RECT 208.910 2574.240 213.830 2574.380 ;
        RECT 208.910 2574.180 209.230 2574.240 ;
        RECT 211.670 2574.180 211.990 2574.240 ;
        RECT 213.510 2574.180 213.830 2574.240 ;
        RECT 210.750 2345.900 211.070 2345.960 ;
        RECT 211.670 2345.900 211.990 2345.960 ;
        RECT 210.750 2345.760 211.990 2345.900 ;
        RECT 210.750 2345.700 211.070 2345.760 ;
        RECT 211.670 2345.700 211.990 2345.760 ;
        RECT 209.830 2221.800 210.150 2221.860 ;
        RECT 211.210 2221.800 211.530 2221.860 ;
        RECT 209.830 2221.660 211.530 2221.800 ;
        RECT 209.830 2221.600 210.150 2221.660 ;
        RECT 211.210 2221.600 211.530 2221.660 ;
        RECT 209.830 2125.580 210.150 2125.640 ;
        RECT 210.750 2125.580 211.070 2125.640 ;
        RECT 209.830 2125.440 211.070 2125.580 ;
        RECT 209.830 2125.380 210.150 2125.440 ;
        RECT 210.750 2125.380 211.070 2125.440 ;
        RECT 210.750 2056.220 211.070 2056.280 ;
        RECT 213.050 2056.220 213.370 2056.280 ;
        RECT 210.750 2056.080 213.370 2056.220 ;
        RECT 210.750 2056.020 211.070 2056.080 ;
        RECT 213.050 2056.020 213.370 2056.080 ;
        RECT 3367.730 2010.660 3368.050 2010.720 ;
        RECT 3376.930 2010.660 3377.250 2010.720 ;
        RECT 3367.730 2010.520 3377.250 2010.660 ;
        RECT 3367.730 2010.460 3368.050 2010.520 ;
        RECT 3376.930 2010.460 3377.250 2010.520 ;
        RECT 208.910 1965.100 209.230 1965.160 ;
        RECT 213.050 1965.100 213.370 1965.160 ;
        RECT 208.910 1964.960 213.370 1965.100 ;
        RECT 208.910 1964.900 209.230 1964.960 ;
        RECT 213.050 1964.900 213.370 1964.960 ;
        RECT 211.670 1960.000 211.990 1960.060 ;
        RECT 213.050 1960.000 213.370 1960.060 ;
        RECT 211.670 1959.860 213.370 1960.000 ;
        RECT 211.670 1959.800 211.990 1959.860 ;
        RECT 213.050 1959.800 213.370 1959.860 ;
        RECT 3367.730 1405.800 3368.050 1405.860 ;
        RECT 3376.930 1405.800 3377.250 1405.860 ;
        RECT 3367.730 1405.660 3377.250 1405.800 ;
        RECT 3367.730 1405.600 3368.050 1405.660 ;
        RECT 3376.930 1405.600 3377.250 1405.660 ;
        RECT 3367.730 794.480 3368.050 794.540 ;
        RECT 3376.470 794.480 3376.790 794.540 ;
        RECT 3367.730 794.340 3376.790 794.480 ;
        RECT 3367.730 794.280 3368.050 794.340 ;
        RECT 3376.470 794.280 3376.790 794.340 ;
        RECT 208.910 748.240 209.230 748.300 ;
        RECT 211.670 748.240 211.990 748.300 ;
        RECT 208.910 748.100 211.990 748.240 ;
        RECT 208.910 748.040 209.230 748.100 ;
        RECT 211.670 748.040 211.990 748.100 ;
        RECT 210.750 704.040 211.070 704.100 ;
        RECT 211.670 704.040 211.990 704.100 ;
        RECT 210.750 703.900 211.990 704.040 ;
        RECT 210.750 703.840 211.070 703.900 ;
        RECT 211.670 703.840 211.990 703.900 ;
        RECT 210.750 676.160 211.070 676.220 ;
        RECT 211.210 676.160 211.530 676.220 ;
        RECT 210.750 676.020 211.530 676.160 ;
        RECT 210.750 675.960 211.070 676.020 ;
        RECT 211.210 675.960 211.530 676.020 ;
        RECT 210.750 579.940 211.070 580.000 ;
        RECT 211.670 579.940 211.990 580.000 ;
        RECT 210.750 579.800 211.990 579.940 ;
        RECT 210.750 579.740 211.070 579.800 ;
        RECT 211.670 579.740 211.990 579.800 ;
        RECT 210.750 482.500 211.070 482.760 ;
        RECT 210.840 482.360 210.980 482.500 ;
        RECT 211.670 482.360 211.990 482.420 ;
        RECT 210.840 482.220 211.990 482.360 ;
        RECT 211.670 482.160 211.990 482.220 ;
        RECT 211.670 317.460 211.990 317.520 ;
        RECT 213.050 317.460 213.370 317.520 ;
        RECT 211.670 317.320 213.370 317.460 ;
        RECT 211.670 317.260 211.990 317.320 ;
        RECT 213.050 317.260 213.370 317.320 ;
        RECT 213.050 228.040 213.370 228.100 ;
        RECT 1271.510 228.040 1271.830 228.100 ;
        RECT 213.050 227.900 1271.830 228.040 ;
        RECT 213.050 227.840 213.370 227.900 ;
        RECT 1271.510 227.840 1271.830 227.900 ;
        RECT 1820.750 227.700 1821.070 227.760 ;
        RECT 3367.730 227.700 3368.050 227.760 ;
        RECT 1820.750 227.560 3368.050 227.700 ;
        RECT 1820.750 227.500 1821.070 227.560 ;
        RECT 3367.730 227.500 3368.050 227.560 ;
        RECT 1271.510 221.580 1271.830 221.640 ;
        RECT 1796.830 221.580 1797.150 221.640 ;
        RECT 1818.450 221.580 1818.770 221.640 ;
        RECT 1820.750 221.580 1821.070 221.640 ;
        RECT 1271.510 221.440 1821.070 221.580 ;
        RECT 1271.510 221.380 1271.830 221.440 ;
        RECT 1796.830 221.380 1797.150 221.440 ;
        RECT 1818.450 221.380 1818.770 221.440 ;
        RECT 1820.750 221.380 1821.070 221.440 ;
      LAYER via ;
        RECT 1226.460 4953.840 1226.720 4954.100 ;
        RECT 1352.500 4953.840 1352.760 4954.100 ;
        RECT 681.360 4953.500 681.620 4953.760 ;
        RECT 1448.640 4953.500 1448.900 4953.760 ;
        RECT 1572.840 4953.840 1573.100 4954.100 ;
        RECT 1573.300 4953.840 1573.560 4954.100 ;
        RECT 1226.460 4952.820 1226.720 4953.080 ;
        RECT 1862.640 4953.160 1862.900 4953.420 ;
        RECT 2316.660 4953.160 2316.920 4953.420 ;
        RECT 2318.040 4953.160 2318.300 4953.420 ;
        RECT 1766.500 4952.820 1766.760 4953.080 ;
        RECT 1766.500 4951.460 1766.760 4951.720 ;
        RECT 1771.560 4951.460 1771.820 4951.720 ;
        RECT 1862.640 4951.460 1862.900 4951.720 ;
        RECT 2318.040 4950.440 2318.300 4950.700 ;
        RECT 3367.300 4950.100 3367.560 4950.360 ;
        RECT 3367.300 3839.320 3367.560 3839.580 ;
        RECT 3376.960 3839.320 3377.220 3839.580 ;
        RECT 208.940 3786.280 209.200 3786.540 ;
        RECT 212.620 3786.280 212.880 3786.540 ;
        RECT 3367.760 3726.440 3368.020 3726.700 ;
        RECT 3376.040 3726.440 3376.300 3726.700 ;
        RECT 213.080 3238.880 213.340 3239.140 ;
        RECT 212.160 3237.520 212.420 3237.780 ;
        RECT 3367.760 3231.400 3368.020 3231.660 ;
        RECT 3376.960 3231.400 3377.220 3231.660 ;
        RECT 212.160 3215.080 212.420 3215.340 ;
        RECT 213.540 3215.080 213.800 3215.340 ;
        RECT 208.940 3178.360 209.200 3178.620 ;
        RECT 211.240 3178.360 211.500 3178.620 ;
        RECT 213.540 3178.360 213.800 3178.620 ;
        RECT 210.780 3091.320 211.040 3091.580 ;
        RECT 211.700 3091.320 211.960 3091.580 ;
        RECT 210.780 3090.640 211.040 3090.900 ;
        RECT 211.700 3090.640 211.960 3090.900 ;
        RECT 210.780 2994.760 211.040 2995.020 ;
        RECT 212.160 2994.760 212.420 2995.020 ;
        RECT 212.160 2897.860 212.420 2898.120 ;
        RECT 213.080 2897.860 213.340 2898.120 ;
        RECT 212.160 2801.300 212.420 2801.560 ;
        RECT 213.540 2801.300 213.800 2801.560 ;
        RECT 213.540 2787.360 213.800 2787.620 ;
        RECT 214.000 2787.360 214.260 2787.620 ;
        RECT 3367.760 2617.700 3368.020 2617.960 ;
        RECT 3376.960 2617.700 3377.220 2617.960 ;
        RECT 208.940 2574.180 209.200 2574.440 ;
        RECT 211.700 2574.180 211.960 2574.440 ;
        RECT 213.540 2574.180 213.800 2574.440 ;
        RECT 210.780 2345.700 211.040 2345.960 ;
        RECT 211.700 2345.700 211.960 2345.960 ;
        RECT 209.860 2221.600 210.120 2221.860 ;
        RECT 211.240 2221.600 211.500 2221.860 ;
        RECT 209.860 2125.380 210.120 2125.640 ;
        RECT 210.780 2125.380 211.040 2125.640 ;
        RECT 210.780 2056.020 211.040 2056.280 ;
        RECT 213.080 2056.020 213.340 2056.280 ;
        RECT 3367.760 2010.460 3368.020 2010.720 ;
        RECT 3376.960 2010.460 3377.220 2010.720 ;
        RECT 208.940 1964.900 209.200 1965.160 ;
        RECT 213.080 1964.900 213.340 1965.160 ;
        RECT 211.700 1959.800 211.960 1960.060 ;
        RECT 213.080 1959.800 213.340 1960.060 ;
        RECT 3367.760 1405.600 3368.020 1405.860 ;
        RECT 3376.960 1405.600 3377.220 1405.860 ;
        RECT 3367.760 794.280 3368.020 794.540 ;
        RECT 3376.500 794.280 3376.760 794.540 ;
        RECT 208.940 748.040 209.200 748.300 ;
        RECT 211.700 748.040 211.960 748.300 ;
        RECT 210.780 703.840 211.040 704.100 ;
        RECT 211.700 703.840 211.960 704.100 ;
        RECT 210.780 675.960 211.040 676.220 ;
        RECT 211.240 675.960 211.500 676.220 ;
        RECT 210.780 579.740 211.040 580.000 ;
        RECT 211.700 579.740 211.960 580.000 ;
        RECT 210.780 482.500 211.040 482.760 ;
        RECT 211.700 482.160 211.960 482.420 ;
        RECT 211.700 317.260 211.960 317.520 ;
        RECT 213.080 317.260 213.340 317.520 ;
        RECT 213.080 227.840 213.340 228.100 ;
        RECT 1271.540 227.840 1271.800 228.100 ;
        RECT 1820.780 227.500 1821.040 227.760 ;
        RECT 3367.760 227.500 3368.020 227.760 ;
        RECT 1271.540 221.380 1271.800 221.640 ;
        RECT 1796.860 221.380 1797.120 221.640 ;
        RECT 1818.480 221.380 1818.740 221.640 ;
        RECT 1820.780 221.380 1821.040 221.640 ;
      LAYER met2 ;
        RECT 681.445 4977.260 681.725 4979.435 ;
        RECT 681.420 4977.035 681.725 4977.260 ;
        RECT 1226.445 4977.035 1226.725 4979.435 ;
        RECT 1771.445 4977.260 1771.725 4979.435 ;
        RECT 2316.445 4977.330 2316.725 4979.435 ;
        RECT 1771.445 4977.035 1771.760 4977.260 ;
        RECT 2316.445 4977.035 2316.860 4977.330 ;
        RECT 681.420 4953.790 681.560 4977.035 ;
        RECT 1226.520 4954.130 1226.660 4977.035 ;
        RECT 1226.460 4953.810 1226.720 4954.130 ;
        RECT 1352.490 4953.955 1352.770 4954.325 ;
        RECT 1448.630 4953.955 1448.910 4954.325 ;
        RECT 1572.900 4954.130 1573.500 4954.210 ;
        RECT 1572.840 4954.070 1573.560 4954.130 ;
        RECT 1352.500 4953.810 1352.760 4953.955 ;
        RECT 681.360 4953.470 681.620 4953.790 ;
        RECT 1226.520 4953.110 1226.660 4953.810 ;
        RECT 1448.700 4953.790 1448.840 4953.955 ;
        RECT 1572.840 4953.810 1573.100 4954.070 ;
        RECT 1573.300 4953.810 1573.560 4954.070 ;
        RECT 1448.640 4953.470 1448.900 4953.790 ;
        RECT 1226.460 4952.790 1226.720 4953.110 ;
        RECT 1766.500 4952.790 1766.760 4953.110 ;
        RECT 1766.560 4951.750 1766.700 4952.790 ;
        RECT 1771.620 4951.750 1771.760 4977.035 ;
        RECT 2316.720 4953.450 2316.860 4977.035 ;
        RECT 1862.640 4953.130 1862.900 4953.450 ;
        RECT 2316.660 4953.130 2316.920 4953.450 ;
        RECT 2318.040 4953.130 2318.300 4953.450 ;
        RECT 1862.700 4951.750 1862.840 4953.130 ;
        RECT 1766.500 4951.430 1766.760 4951.750 ;
        RECT 1771.560 4951.430 1771.820 4951.750 ;
        RECT 1862.640 4951.430 1862.900 4951.750 ;
        RECT 2318.100 4950.730 2318.240 4953.130 ;
        RECT 2318.040 4950.410 2318.300 4950.730 ;
        RECT 3367.300 4950.070 3367.560 4950.390 ;
        RECT 3367.360 3839.610 3367.500 4950.070 ;
        RECT 3367.300 3839.290 3367.560 3839.610 ;
        RECT 3376.960 3839.290 3377.220 3839.610 ;
        RECT 3377.020 3837.555 3377.160 3839.290 ;
        RECT 3377.020 3837.485 3379.435 3837.555 ;
        RECT 3376.100 3837.345 3379.435 3837.485 ;
        RECT 208.565 3788.445 210.965 3788.725 ;
        RECT 209.000 3786.570 209.140 3788.445 ;
        RECT 208.940 3786.250 209.200 3786.570 ;
        RECT 212.620 3786.250 212.880 3786.570 ;
        RECT 212.680 3312.010 212.820 3786.250 ;
        RECT 3376.100 3726.730 3376.240 3837.345 ;
        RECT 3377.035 3837.275 3379.435 3837.345 ;
        RECT 3367.760 3726.410 3368.020 3726.730 ;
        RECT 3376.040 3726.410 3376.300 3726.730 ;
        RECT 212.680 3311.870 213.280 3312.010 ;
        RECT 213.140 3239.170 213.280 3311.870 ;
        RECT 213.080 3238.850 213.340 3239.170 ;
        RECT 212.160 3237.490 212.420 3237.810 ;
        RECT 212.220 3215.370 212.360 3237.490 ;
        RECT 3367.820 3231.690 3367.960 3726.410 ;
        RECT 3367.760 3231.370 3368.020 3231.690 ;
        RECT 3376.960 3231.370 3377.220 3231.690 ;
        RECT 212.160 3215.050 212.420 3215.370 ;
        RECT 213.540 3215.050 213.800 3215.370 ;
        RECT 208.610 3180.725 209.140 3180.770 ;
        RECT 208.565 3180.445 210.965 3180.725 ;
        RECT 209.000 3178.650 209.140 3180.445 ;
        RECT 213.600 3178.650 213.740 3215.050 ;
        RECT 208.940 3178.330 209.200 3178.650 ;
        RECT 211.240 3178.330 211.500 3178.650 ;
        RECT 213.540 3178.330 213.800 3178.650 ;
        RECT 211.300 3167.850 211.440 3178.330 ;
        RECT 210.840 3167.710 211.440 3167.850 ;
        RECT 210.840 3091.610 210.980 3167.710 ;
        RECT 210.780 3091.290 211.040 3091.610 ;
        RECT 211.700 3091.290 211.960 3091.610 ;
        RECT 211.760 3090.930 211.900 3091.290 ;
        RECT 210.780 3090.610 211.040 3090.930 ;
        RECT 211.700 3090.610 211.960 3090.930 ;
        RECT 210.840 2995.050 210.980 3090.610 ;
        RECT 210.780 2994.730 211.040 2995.050 ;
        RECT 212.160 2994.730 212.420 2995.050 ;
        RECT 212.220 2925.770 212.360 2994.730 ;
        RECT 212.220 2925.630 213.280 2925.770 ;
        RECT 213.140 2898.150 213.280 2925.630 ;
        RECT 212.160 2897.830 212.420 2898.150 ;
        RECT 213.080 2897.830 213.340 2898.150 ;
        RECT 212.220 2801.590 212.360 2897.830 ;
        RECT 212.160 2801.270 212.420 2801.590 ;
        RECT 213.540 2801.270 213.800 2801.590 ;
        RECT 213.600 2787.650 213.740 2801.270 ;
        RECT 213.540 2787.330 213.800 2787.650 ;
        RECT 214.000 2787.330 214.260 2787.650 ;
        RECT 214.060 2691.170 214.200 2787.330 ;
        RECT 214.060 2691.030 214.660 2691.170 ;
        RECT 214.520 2636.090 214.660 2691.030 ;
        RECT 213.600 2635.950 214.660 2636.090 ;
        RECT 213.600 2574.470 213.740 2635.950 ;
        RECT 3367.820 2617.990 3367.960 3231.370 ;
        RECT 3377.020 3229.555 3377.160 3231.370 ;
        RECT 3377.020 3229.415 3379.435 3229.555 ;
        RECT 3377.035 3229.275 3379.435 3229.415 ;
        RECT 3377.035 2620.380 3379.435 2620.555 ;
        RECT 3377.020 2620.275 3379.435 2620.380 ;
        RECT 3377.020 2617.990 3377.160 2620.275 ;
        RECT 3367.760 2617.670 3368.020 2617.990 ;
        RECT 3376.960 2617.670 3377.220 2617.990 ;
        RECT 208.940 2574.150 209.200 2574.470 ;
        RECT 211.700 2574.150 211.960 2574.470 ;
        RECT 213.540 2574.150 213.800 2574.470 ;
        RECT 209.000 2571.725 209.140 2574.150 ;
        RECT 208.565 2571.445 210.965 2571.725 ;
        RECT 211.760 2483.770 211.900 2574.150 ;
        RECT 211.300 2483.630 211.900 2483.770 ;
        RECT 211.300 2387.890 211.440 2483.630 ;
        RECT 210.840 2387.750 211.440 2387.890 ;
        RECT 210.840 2345.990 210.980 2387.750 ;
        RECT 210.780 2345.670 211.040 2345.990 ;
        RECT 211.700 2345.670 211.960 2345.990 ;
        RECT 211.760 2249.170 211.900 2345.670 ;
        RECT 211.300 2249.030 211.900 2249.170 ;
        RECT 211.300 2221.890 211.440 2249.030 ;
        RECT 209.860 2221.570 210.120 2221.890 ;
        RECT 211.240 2221.570 211.500 2221.890 ;
        RECT 209.920 2125.670 210.060 2221.570 ;
        RECT 209.860 2125.350 210.120 2125.670 ;
        RECT 210.780 2125.350 211.040 2125.670 ;
        RECT 210.840 2056.310 210.980 2125.350 ;
        RECT 210.780 2055.990 211.040 2056.310 ;
        RECT 213.080 2055.990 213.340 2056.310 ;
        RECT 213.140 1965.190 213.280 2055.990 ;
        RECT 3367.820 2010.750 3367.960 2617.670 ;
        RECT 3377.035 2011.415 3379.435 2011.555 ;
        RECT 3377.020 2011.275 3379.435 2011.415 ;
        RECT 3377.020 2010.750 3377.160 2011.275 ;
        RECT 3367.760 2010.430 3368.020 2010.750 ;
        RECT 3376.960 2010.430 3377.220 2010.750 ;
        RECT 208.940 1964.870 209.200 1965.190 ;
        RECT 213.080 1964.870 213.340 1965.190 ;
        RECT 209.000 1962.725 209.140 1964.870 ;
        RECT 208.565 1962.445 210.965 1962.725 ;
        RECT 213.140 1960.090 213.280 1964.870 ;
        RECT 211.700 1959.770 211.960 1960.090 ;
        RECT 213.080 1959.770 213.340 1960.090 ;
        RECT 211.760 1357.010 211.900 1959.770 ;
        RECT 3367.820 1405.890 3367.960 2010.430 ;
        RECT 3367.760 1405.570 3368.020 1405.890 ;
        RECT 3376.960 1405.570 3377.220 1405.890 ;
        RECT 209.000 1356.870 211.900 1357.010 ;
        RECT 209.000 1354.725 209.140 1356.870 ;
        RECT 208.565 1354.445 210.965 1354.725 ;
        RECT 211.760 748.330 211.900 1356.870 ;
        RECT 3367.820 794.570 3367.960 1405.570 ;
        RECT 3377.020 1403.555 3377.160 1405.570 ;
        RECT 3377.020 1403.415 3379.435 1403.555 ;
        RECT 3377.035 1403.275 3379.435 1403.415 ;
        RECT 3367.760 794.250 3368.020 794.570 ;
        RECT 3376.500 794.485 3376.760 794.570 ;
        RECT 3377.035 794.485 3379.435 794.555 ;
        RECT 3376.500 794.345 3379.435 794.485 ;
        RECT 3376.500 794.250 3376.760 794.345 ;
        RECT 3377.035 794.275 3379.435 794.345 ;
        RECT 208.940 748.010 209.200 748.330 ;
        RECT 211.700 748.010 211.960 748.330 ;
        RECT 209.000 745.725 209.140 748.010 ;
        RECT 208.565 745.445 210.965 745.725 ;
        RECT 211.760 704.130 211.900 748.010 ;
        RECT 210.780 703.810 211.040 704.130 ;
        RECT 211.700 703.810 211.960 704.130 ;
        RECT 210.840 703.530 210.980 703.810 ;
        RECT 210.840 703.390 211.440 703.530 ;
        RECT 211.300 676.250 211.440 703.390 ;
        RECT 210.780 675.930 211.040 676.250 ;
        RECT 211.240 675.930 211.500 676.250 ;
        RECT 210.840 580.030 210.980 675.930 ;
        RECT 210.780 579.710 211.040 580.030 ;
        RECT 211.700 579.710 211.960 580.030 ;
        RECT 211.760 531.490 211.900 579.710 ;
        RECT 210.380 531.350 211.900 531.490 ;
        RECT 210.380 483.210 210.520 531.350 ;
        RECT 210.380 483.070 210.980 483.210 ;
        RECT 210.840 482.790 210.980 483.070 ;
        RECT 210.780 482.470 211.040 482.790 ;
        RECT 211.700 482.130 211.960 482.450 ;
        RECT 211.760 317.550 211.900 482.130 ;
        RECT 211.700 317.230 211.960 317.550 ;
        RECT 213.080 317.230 213.340 317.550 ;
        RECT 213.140 228.130 213.280 317.230 ;
        RECT 213.080 227.810 213.340 228.130 ;
        RECT 1271.540 227.810 1271.800 228.130 ;
        RECT 1271.600 221.670 1271.740 227.810 ;
        RECT 3367.820 227.790 3367.960 794.250 ;
        RECT 1820.780 227.470 1821.040 227.790 ;
        RECT 3367.760 227.470 3368.020 227.790 ;
        RECT 1820.840 221.670 1820.980 227.470 ;
        RECT 1271.540 221.350 1271.800 221.670 ;
        RECT 1796.860 221.350 1797.120 221.670 ;
        RECT 1818.480 221.350 1818.740 221.670 ;
        RECT 1820.780 221.350 1821.040 221.670 ;
        RECT 1271.600 201.010 1271.740 221.350 ;
        RECT 1796.920 210.965 1797.060 221.350 ;
        RECT 1818.540 210.965 1818.680 221.350 ;
        RECT 1796.655 209.030 1797.060 210.965 ;
        RECT 1818.275 209.030 1818.680 210.965 ;
        RECT 1796.655 208.565 1796.935 209.030 ;
        RECT 1818.275 208.565 1818.555 209.030 ;
        RECT 1271.515 200.870 1271.740 201.010 ;
        RECT 1271.515 200.000 1271.655 200.870 ;
        RECT 1271.455 198.530 1271.715 200.000 ;
      LAYER via2 ;
        RECT 1352.490 4954.000 1352.770 4954.280 ;
        RECT 1448.630 4954.000 1448.910 4954.280 ;
      LAYER met3 ;
        RECT 1352.465 4954.290 1352.795 4954.305 ;
        RECT 1448.605 4954.290 1448.935 4954.305 ;
        RECT 1352.465 4953.990 1448.935 4954.290 ;
        RECT 1352.465 4953.975 1352.795 4953.990 ;
        RECT 1448.605 4953.975 1448.935 4953.990 ;
    END
  END porb_h
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1215.200 33.375 1277.900 95.990 ;
    END
  END resetb
  PIN resetb_core_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1254.335 190.155 1255.065 200.000 ;
        RECT 1254.335 189.855 1255.365 190.155 ;
        RECT 1254.335 189.555 1255.100 189.855 ;
        RECT 1255.365 189.555 1255.830 189.855 ;
        RECT 1254.335 189.090 1255.830 189.555 ;
        RECT 1255.100 185.230 1255.830 189.090 ;
    END
  END resetb_core_h
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3490.140 4389.045 3557.570 4445.685 ;
    END
  END vccd
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2847.200 33.375 2909.900 95.990 ;
    END
  END vdda
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 33.375 4390.100 95.990 4452.800 ;
    END
  END vddio
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 673.200 33.375 735.900 95.990 ;
    END
  END vssa
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2308.045 30.430 2364.685 97.860 ;
    END
  END vssd
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2854.100 5092.010 2916.800 5154.625 ;
    END
  END vssio
  OBS
      LAYER li1 ;
        RECT 667.840 4988.230 748.160 5187.705 ;
        RECT 1212.840 4988.230 1293.160 5187.705 ;
        RECT 1757.840 4988.230 1838.160 5187.705 ;
        RECT 2302.840 4988.230 2383.160 5187.705 ;
        RECT 2849.070 4990.035 2920.775 5187.695 ;
        RECT 0.305 4384.610 197.965 4456.855 ;
        RECT 3391.020 4380.245 3587.780 4454.760 ;
        RECT 0.295 3774.840 199.770 3855.160 ;
        RECT 3388.230 3770.840 3587.705 3851.160 ;
        RECT 0.295 3166.840 199.770 3247.160 ;
        RECT 3388.230 3162.840 3587.705 3243.160 ;
        RECT 0.295 2557.840 199.770 2638.160 ;
        RECT 3388.230 2553.840 3587.705 2634.160 ;
        RECT 0.295 1948.840 199.770 2029.160 ;
        RECT 3388.230 1944.840 3587.705 2025.160 ;
        RECT 0.295 1340.840 199.770 1421.160 ;
        RECT 3388.230 1336.840 3587.705 1417.160 ;
        RECT 0.295 731.840 199.770 812.160 ;
        RECT 3388.230 727.840 3587.705 808.160 ;
        RECT 669.225 0.305 740.930 197.965 ;
        RECT 1209.000 0.780 1284.000 199.815 ;
        RECT 1751.840 0.295 1832.160 199.770 ;
        RECT 2299.245 0.220 2373.760 196.980 ;
        RECT 2843.145 0.305 2915.390 197.965 ;
      LAYER met1 ;
        RECT 667.855 4981.155 748.145 5188.000 ;
        RECT 1212.855 4981.155 1293.145 5188.000 ;
        RECT 1757.855 4981.155 1838.145 5188.000 ;
        RECT 2302.855 4981.155 2383.145 5188.000 ;
        RECT 2848.185 4990.035 2921.620 5187.725 ;
      LAYER met1 ;
        RECT 707.090 4978.180 707.410 4978.240 ;
        RECT 745.730 4978.180 746.050 4978.240 ;
        RECT 707.090 4978.040 746.050 4978.180 ;
        RECT 707.090 4977.980 707.410 4978.040 ;
        RECT 745.730 4977.980 746.050 4978.040 ;
        RECT 2341.930 4977.500 2342.250 4977.560 ;
        RECT 2380.570 4977.500 2380.890 4977.560 ;
        RECT 2341.930 4977.360 2380.890 4977.500 ;
        RECT 2341.930 4977.300 2342.250 4977.360 ;
        RECT 2380.570 4977.300 2380.890 4977.360 ;
        RECT 1251.730 4977.160 1252.050 4977.220 ;
        RECT 1290.830 4977.160 1291.150 4977.220 ;
        RECT 1251.730 4977.020 1291.150 4977.160 ;
        RECT 1251.730 4976.960 1252.050 4977.020 ;
        RECT 1290.830 4976.960 1291.150 4977.020 ;
        RECT 1228.270 4960.500 1228.590 4960.560 ;
        RECT 1282.090 4960.500 1282.410 4960.560 ;
        RECT 1228.270 4960.360 1282.410 4960.500 ;
        RECT 1228.270 4960.300 1228.590 4960.360 ;
        RECT 1282.090 4960.300 1282.410 4960.360 ;
        RECT 684.550 4954.040 684.870 4954.100 ;
        RECT 1225.970 4954.040 1226.290 4954.100 ;
        RECT 684.550 4953.900 1226.290 4954.040 ;
        RECT 684.550 4953.840 684.870 4953.900 ;
        RECT 1225.970 4953.840 1226.290 4953.900 ;
        RECT 1796.370 4954.040 1796.690 4954.100 ;
        RECT 1836.390 4954.040 1836.710 4954.100 ;
        RECT 2369.990 4954.040 2370.310 4954.100 ;
        RECT 2372.290 4954.040 2372.610 4954.100 ;
        RECT 1796.370 4953.900 1836.710 4954.040 ;
        RECT 1796.370 4953.840 1796.690 4953.900 ;
        RECT 1836.390 4953.840 1836.710 4953.900 ;
        RECT 1836.940 4953.900 2372.610 4954.040 ;
        RECT 1827.190 4953.700 1827.510 4953.760 ;
        RECT 1836.940 4953.700 1837.080 4953.900 ;
        RECT 2369.990 4953.840 2370.310 4953.900 ;
        RECT 2372.290 4953.840 2372.610 4953.900 ;
        RECT 2319.850 4953.700 2320.170 4953.760 ;
        RECT 2856.670 4953.700 2856.990 4953.760 ;
        RECT 1827.190 4953.560 1837.080 4953.700 ;
        RECT 1837.400 4953.560 2856.990 4953.700 ;
        RECT 1827.190 4953.500 1827.510 4953.560 ;
        RECT 1089.810 4953.360 1090.130 4953.420 ;
        RECT 993.300 4953.220 1090.130 4953.360 ;
        RECT 993.300 4953.020 993.440 4953.220 ;
        RECT 1089.810 4953.160 1090.130 4953.220 ;
        RECT 897.160 4952.880 993.440 4953.020 ;
        RECT 662.470 4952.680 662.790 4952.740 ;
        RECT 623.920 4952.540 662.790 4952.680 ;
        RECT 224.090 4952.340 224.410 4952.400 ;
        RECT 317.470 4952.340 317.790 4952.400 ;
        RECT 224.090 4952.200 317.790 4952.340 ;
        RECT 224.090 4952.140 224.410 4952.200 ;
        RECT 317.470 4952.140 317.790 4952.200 ;
        RECT 412.230 4952.340 412.550 4952.400 ;
        RECT 623.920 4952.340 624.060 4952.540 ;
        RECT 662.470 4952.480 662.790 4952.540 ;
        RECT 736.990 4952.680 737.310 4952.740 ;
        RECT 897.160 4952.680 897.300 4952.880 ;
        RECT 736.990 4952.540 897.300 4952.680 ;
        RECT 1282.090 4952.680 1282.410 4952.740 ;
        RECT 1435.270 4952.680 1435.590 4952.740 ;
        RECT 1282.090 4952.540 1435.590 4952.680 ;
        RECT 736.990 4952.480 737.310 4952.540 ;
        RECT 1282.090 4952.480 1282.410 4952.540 ;
        RECT 1435.270 4952.480 1435.590 4952.540 ;
        RECT 1545.210 4952.680 1545.530 4952.740 ;
        RECT 1628.470 4952.680 1628.790 4952.740 ;
        RECT 1545.210 4952.540 1628.790 4952.680 ;
        RECT 1545.210 4952.480 1545.530 4952.540 ;
        RECT 1628.470 4952.480 1628.790 4952.540 ;
        RECT 1738.410 4952.680 1738.730 4952.740 ;
        RECT 1827.190 4952.680 1827.510 4952.740 ;
        RECT 1738.410 4952.540 1827.510 4952.680 ;
        RECT 1738.410 4952.480 1738.730 4952.540 ;
        RECT 1827.190 4952.480 1827.510 4952.540 ;
        RECT 412.230 4952.200 510.900 4952.340 ;
        RECT 412.230 4952.140 412.550 4952.200 ;
        RECT 224.550 4951.660 224.870 4951.720 ;
        RECT 224.550 4951.520 318.620 4951.660 ;
        RECT 224.550 4951.460 224.870 4951.520 ;
        RECT 318.480 4951.320 318.620 4951.520 ;
        RECT 386.470 4951.320 386.790 4951.380 ;
        RECT 510.760 4951.320 510.900 4952.200 ;
        RECT 565.960 4952.200 624.060 4952.340 ;
        RECT 530.910 4952.000 531.230 4952.060 ;
        RECT 565.960 4952.000 566.100 4952.200 ;
        RECT 772.870 4952.140 773.190 4952.400 ;
        RECT 1225.970 4952.340 1226.290 4952.400 ;
        RECT 1229.650 4952.340 1229.970 4952.400 ;
        RECT 1448.610 4952.340 1448.930 4952.400 ;
        RECT 1225.970 4952.200 1448.930 4952.340 ;
        RECT 1225.970 4952.140 1226.290 4952.200 ;
        RECT 1229.650 4952.140 1229.970 4952.200 ;
        RECT 1448.610 4952.140 1448.930 4952.200 ;
        RECT 1449.530 4952.340 1449.850 4952.400 ;
        RECT 1774.750 4952.340 1775.070 4952.400 ;
        RECT 1837.400 4952.340 1837.540 4953.560 ;
        RECT 2319.850 4953.500 2320.170 4953.560 ;
        RECT 2856.670 4953.500 2856.990 4953.560 ;
        RECT 1449.530 4952.200 1837.540 4952.340 ;
        RECT 1449.530 4952.140 1449.850 4952.200 ;
        RECT 1774.750 4952.140 1775.070 4952.200 ;
        RECT 530.910 4951.860 566.100 4952.000 ;
        RECT 758.610 4952.000 758.930 4952.060 ;
        RECT 772.960 4952.000 773.100 4952.140 ;
        RECT 758.610 4951.860 773.100 4952.000 ;
        RECT 1179.510 4952.000 1179.830 4952.060 ;
        RECT 1227.810 4952.000 1228.130 4952.060 ;
        RECT 1179.510 4951.860 1228.130 4952.000 ;
        RECT 530.910 4951.800 531.230 4951.860 ;
        RECT 758.610 4951.800 758.930 4951.860 ;
        RECT 1179.510 4951.800 1179.830 4951.860 ;
        RECT 1227.810 4951.800 1228.130 4951.860 ;
        RECT 1449.990 4952.000 1450.310 4952.060 ;
        RECT 1545.210 4952.000 1545.530 4952.060 ;
        RECT 1449.990 4951.860 1545.530 4952.000 ;
        RECT 1449.990 4951.800 1450.310 4951.860 ;
        RECT 1545.210 4951.800 1545.530 4951.860 ;
        RECT 662.930 4951.320 663.250 4951.380 ;
        RECT 758.610 4951.320 758.930 4951.380 ;
        RECT 966.070 4951.320 966.390 4951.380 ;
        RECT 318.480 4951.180 386.790 4951.320 ;
        RECT 386.470 4951.120 386.790 4951.180 ;
        RECT 412.780 4951.180 435.000 4951.320 ;
        RECT 510.760 4951.180 607.040 4951.320 ;
        RECT 317.470 4950.980 317.790 4951.040 ;
        RECT 412.230 4950.980 412.550 4951.040 ;
        RECT 317.470 4950.840 412.550 4950.980 ;
        RECT 317.470 4950.780 317.790 4950.840 ;
        RECT 412.230 4950.780 412.550 4950.840 ;
        RECT 211.210 4950.640 211.530 4950.700 ;
        RECT 412.780 4950.640 412.920 4951.180 ;
        RECT 211.210 4950.500 412.920 4950.640 ;
        RECT 211.210 4950.440 211.530 4950.500 ;
        RECT 414.070 4950.440 414.390 4950.700 ;
        RECT 434.860 4950.640 435.000 4951.180 ;
        RECT 606.900 4950.980 607.040 4951.180 ;
        RECT 662.930 4951.180 758.930 4951.320 ;
        RECT 662.930 4951.120 663.250 4951.180 ;
        RECT 758.610 4951.120 758.930 4951.180 ;
        RECT 896.700 4951.180 966.390 4951.320 ;
        RECT 684.550 4950.980 684.870 4951.040 ;
        RECT 606.900 4950.840 684.870 4950.980 ;
        RECT 684.550 4950.780 684.870 4950.840 ;
        RECT 773.330 4950.980 773.650 4951.040 ;
        RECT 773.330 4950.840 869.240 4950.980 ;
        RECT 773.330 4950.780 773.650 4950.840 ;
        RECT 510.670 4950.640 510.990 4950.700 ;
        RECT 434.860 4950.500 510.990 4950.640 ;
        RECT 510.670 4950.440 510.990 4950.500 ;
        RECT 530.910 4950.440 531.230 4950.700 ;
        RECT 531.370 4950.640 531.690 4950.700 ;
        RECT 736.990 4950.640 737.310 4950.700 ;
        RECT 531.370 4950.500 737.310 4950.640 ;
        RECT 869.100 4950.640 869.240 4950.840 ;
        RECT 896.700 4950.640 896.840 4951.180 ;
        RECT 966.070 4951.120 966.390 4951.180 ;
        RECT 1089.810 4951.320 1090.130 4951.380 ;
        RECT 1227.350 4951.320 1227.670 4951.380 ;
        RECT 1228.270 4951.320 1228.590 4951.380 ;
        RECT 1089.810 4951.180 1179.740 4951.320 ;
        RECT 1089.810 4951.120 1090.130 4951.180 ;
        RECT 1179.600 4950.980 1179.740 4951.180 ;
        RECT 1227.350 4951.180 1228.590 4951.320 ;
        RECT 1227.350 4951.120 1227.670 4951.180 ;
        RECT 1228.270 4951.120 1228.590 4951.180 ;
        RECT 1380.070 4951.320 1380.390 4951.380 ;
        RECT 1474.830 4951.320 1475.150 4951.380 ;
        RECT 1380.070 4951.180 1475.150 4951.320 ;
        RECT 1380.070 4951.120 1380.390 4951.180 ;
        RECT 1474.830 4951.120 1475.150 4951.180 ;
        RECT 1226.890 4950.980 1227.210 4951.040 ;
        RECT 1179.600 4950.840 1227.210 4950.980 ;
        RECT 1226.890 4950.780 1227.210 4950.840 ;
        RECT 1227.810 4950.980 1228.130 4951.040 ;
        RECT 1379.610 4950.980 1379.930 4951.040 ;
        RECT 1227.810 4950.840 1379.930 4950.980 ;
        RECT 1227.810 4950.780 1228.130 4950.840 ;
        RECT 1379.610 4950.780 1379.930 4950.840 ;
        RECT 2856.670 4950.980 2856.990 4951.040 ;
        RECT 2870.010 4950.980 2870.330 4951.040 ;
        RECT 3373.710 4950.980 3374.030 4951.040 ;
        RECT 2856.670 4950.840 3374.030 4950.980 ;
        RECT 2856.670 4950.780 2856.990 4950.840 ;
        RECT 2870.010 4950.780 2870.330 4950.840 ;
        RECT 3373.710 4950.780 3374.030 4950.840 ;
        RECT 869.100 4950.500 896.840 4950.640 ;
        RECT 1091.190 4950.640 1091.510 4950.700 ;
        RECT 1179.510 4950.640 1179.830 4950.700 ;
        RECT 1091.190 4950.500 1179.830 4950.640 ;
        RECT 531.370 4950.440 531.690 4950.500 ;
        RECT 736.990 4950.440 737.310 4950.500 ;
        RECT 1091.190 4950.440 1091.510 4950.500 ;
        RECT 1179.510 4950.440 1179.830 4950.500 ;
        RECT 2369.990 4950.640 2370.310 4950.700 ;
        RECT 3365.430 4950.640 3365.750 4950.700 ;
        RECT 2369.990 4950.500 3365.750 4950.640 ;
        RECT 2369.990 4950.440 2370.310 4950.500 ;
        RECT 3365.430 4950.440 3365.750 4950.500 ;
        RECT 414.160 4950.300 414.300 4950.440 ;
        RECT 531.000 4950.300 531.140 4950.440 ;
        RECT 414.160 4950.160 531.140 4950.300 ;
        RECT 222.250 4574.600 222.570 4574.660 ;
        RECT 224.090 4574.600 224.410 4574.660 ;
        RECT 222.250 4574.460 224.410 4574.600 ;
        RECT 222.250 4574.400 222.570 4574.460 ;
        RECT 224.090 4574.400 224.410 4574.460 ;
        RECT 3368.650 4471.580 3368.970 4471.640 ;
        RECT 3373.710 4471.580 3374.030 4471.640 ;
        RECT 3390.270 4471.580 3390.590 4471.640 ;
        RECT 3368.650 4471.440 3390.590 4471.580 ;
        RECT 3368.650 4471.380 3368.970 4471.440 ;
        RECT 3373.710 4471.380 3374.030 4471.440 ;
        RECT 3390.270 4471.380 3390.590 4471.440 ;
      LAYER met1 ;
        RECT 0.275 4384.185 197.965 4456.915 ;
      LAYER met1 ;
        RECT 222.250 4443.700 222.570 4443.760 ;
        RECT 223.630 4443.700 223.950 4443.760 ;
        RECT 222.250 4443.560 223.950 4443.700 ;
        RECT 222.250 4443.500 222.570 4443.560 ;
        RECT 223.630 4443.500 223.950 4443.560 ;
        RECT 3365.430 4400.180 3365.750 4400.240 ;
        RECT 3368.190 4400.180 3368.510 4400.240 ;
        RECT 3365.430 4400.040 3368.510 4400.180 ;
        RECT 3365.430 4399.980 3365.750 4400.040 ;
        RECT 3368.190 4399.980 3368.510 4400.040 ;
        RECT 3368.190 4380.800 3368.510 4380.860 ;
        RECT 3389.350 4380.800 3389.670 4380.860 ;
        RECT 3368.190 4380.660 3389.670 4380.800 ;
        RECT 3368.190 4380.600 3368.510 4380.660 ;
        RECT 3389.350 4380.600 3389.670 4380.660 ;
      LAYER met1 ;
        RECT 3390.035 4380.215 3587.840 4454.880 ;
      LAYER met1 ;
        RECT 3373.710 4374.680 3374.030 4374.740 ;
        RECT 3388.430 4374.680 3388.750 4374.740 ;
        RECT 3373.710 4374.540 3388.750 4374.680 ;
        RECT 3373.710 4374.480 3374.030 4374.540 ;
        RECT 3388.430 4374.480 3388.750 4374.540 ;
        RECT 210.750 4347.140 211.070 4347.200 ;
        RECT 223.630 4347.140 223.950 4347.200 ;
        RECT 210.750 4347.000 223.950 4347.140 ;
        RECT 210.750 4346.940 211.070 4347.000 ;
        RECT 223.630 4346.940 223.950 4347.000 ;
        RECT 223.630 4181.560 223.950 4181.620 ;
        RECT 223.260 4181.420 223.950 4181.560 ;
        RECT 223.260 4181.280 223.400 4181.420 ;
        RECT 223.630 4181.360 223.950 4181.420 ;
        RECT 223.170 4181.020 223.490 4181.280 ;
        RECT 223.170 4154.020 223.490 4154.080 ;
        RECT 223.630 4154.020 223.950 4154.080 ;
        RECT 223.170 4153.880 223.950 4154.020 ;
        RECT 223.170 4153.820 223.490 4153.880 ;
        RECT 223.630 4153.820 223.950 4153.880 ;
        RECT 222.250 3891.680 222.570 3891.940 ;
        RECT 222.340 3891.200 222.480 3891.680 ;
        RECT 222.710 3891.200 223.030 3891.260 ;
        RECT 222.340 3891.060 223.030 3891.200 ;
        RECT 222.710 3891.000 223.030 3891.060 ;
        RECT 211.210 3871.480 211.530 3871.540 ;
        RECT 212.590 3871.480 212.910 3871.540 ;
        RECT 211.210 3871.340 212.910 3871.480 ;
        RECT 211.210 3871.280 211.530 3871.340 ;
        RECT 212.590 3871.280 212.910 3871.340 ;
      LAYER met1 ;
        RECT 0.000 3774.855 206.845 3855.145 ;
      LAYER met1 ;
        RECT 208.910 3846.320 209.230 3846.380 ;
        RECT 212.590 3846.320 212.910 3846.380 ;
        RECT 208.910 3846.180 212.910 3846.320 ;
        RECT 208.910 3846.120 209.230 3846.180 ;
        RECT 212.590 3846.120 212.910 3846.180 ;
        RECT 211.670 3836.800 211.990 3836.860 ;
        RECT 212.590 3836.800 212.910 3836.860 ;
        RECT 211.670 3836.660 212.910 3836.800 ;
        RECT 211.670 3836.600 211.990 3836.660 ;
        RECT 212.590 3836.600 212.910 3836.660 ;
        RECT 3368.650 3836.800 3368.970 3836.860 ;
        RECT 3376.930 3836.800 3377.250 3836.860 ;
        RECT 3368.650 3836.660 3377.250 3836.800 ;
        RECT 3368.650 3836.600 3368.970 3836.660 ;
        RECT 3376.930 3836.600 3377.250 3836.660 ;
        RECT 208.910 3792.600 209.230 3792.660 ;
        RECT 213.050 3792.600 213.370 3792.660 ;
        RECT 220.870 3792.600 221.190 3792.660 ;
        RECT 208.910 3792.460 221.190 3792.600 ;
        RECT 208.910 3792.400 209.230 3792.460 ;
        RECT 213.050 3792.400 213.370 3792.460 ;
        RECT 220.870 3792.400 221.190 3792.460 ;
        RECT 3367.270 3779.680 3367.590 3779.740 ;
        RECT 3368.190 3779.680 3368.510 3779.740 ;
        RECT 3376.930 3779.680 3377.250 3779.740 ;
        RECT 3367.270 3779.540 3377.250 3779.680 ;
        RECT 3367.270 3779.480 3367.590 3779.540 ;
        RECT 3368.190 3779.480 3368.510 3779.540 ;
        RECT 3376.930 3779.480 3377.250 3779.540 ;
      LAYER met1 ;
        RECT 3381.155 3770.855 3588.000 3851.145 ;
      LAYER met1 ;
        RECT 211.670 3757.920 211.990 3757.980 ;
        RECT 213.050 3757.920 213.370 3757.980 ;
        RECT 211.670 3757.780 213.370 3757.920 ;
        RECT 211.670 3757.720 211.990 3757.780 ;
        RECT 213.050 3757.720 213.370 3757.780 ;
        RECT 223.630 3698.560 223.950 3698.820 ;
        RECT 223.720 3698.080 223.860 3698.560 ;
        RECT 224.090 3698.080 224.410 3698.140 ;
        RECT 223.720 3697.940 224.410 3698.080 ;
        RECT 224.090 3697.880 224.410 3697.940 ;
        RECT 223.170 3670.540 223.490 3670.600 ;
        RECT 224.090 3670.540 224.410 3670.600 ;
        RECT 223.170 3670.400 224.410 3670.540 ;
        RECT 223.170 3670.340 223.490 3670.400 ;
        RECT 224.090 3670.340 224.410 3670.400 ;
        RECT 223.170 3601.860 223.490 3601.920 ;
        RECT 224.090 3601.860 224.410 3601.920 ;
        RECT 223.170 3601.720 224.410 3601.860 ;
        RECT 223.170 3601.660 223.490 3601.720 ;
        RECT 224.090 3601.660 224.410 3601.720 ;
        RECT 224.090 3505.100 224.410 3505.360 ;
        RECT 224.180 3504.680 224.320 3505.100 ;
        RECT 224.090 3504.420 224.410 3504.680 ;
        RECT 222.250 3463.820 222.570 3463.880 ;
        RECT 224.090 3463.820 224.410 3463.880 ;
        RECT 222.250 3463.680 224.410 3463.820 ;
        RECT 222.250 3463.620 222.570 3463.680 ;
        RECT 224.090 3463.620 224.410 3463.680 ;
        RECT 222.250 3367.600 222.570 3367.660 ;
        RECT 223.630 3367.600 223.950 3367.660 ;
        RECT 222.250 3367.460 223.950 3367.600 ;
        RECT 222.250 3367.400 222.570 3367.460 ;
        RECT 223.630 3367.400 223.950 3367.460 ;
        RECT 223.630 3312.520 223.950 3312.580 ;
        RECT 223.260 3312.380 223.950 3312.520 ;
        RECT 223.260 3311.900 223.400 3312.380 ;
        RECT 223.630 3312.320 223.950 3312.380 ;
        RECT 223.170 3311.640 223.490 3311.900 ;
        RECT 211.210 3254.720 211.530 3254.780 ;
        RECT 212.130 3254.720 212.450 3254.780 ;
        RECT 211.210 3254.580 212.450 3254.720 ;
        RECT 211.210 3254.520 211.530 3254.580 ;
        RECT 212.130 3254.520 212.450 3254.580 ;
      LAYER met1 ;
        RECT 0.000 3166.855 206.845 3247.145 ;
      LAYER met1 ;
        RECT 208.910 3238.400 209.230 3238.460 ;
        RECT 212.130 3238.400 212.450 3238.460 ;
        RECT 213.050 3238.400 213.370 3238.460 ;
        RECT 208.910 3238.260 213.370 3238.400 ;
        RECT 208.910 3238.200 209.230 3238.260 ;
        RECT 212.130 3238.200 212.450 3238.260 ;
        RECT 213.050 3238.200 213.370 3238.260 ;
        RECT 3368.650 3228.880 3368.970 3228.940 ;
        RECT 3376.930 3228.880 3377.250 3228.940 ;
        RECT 3368.650 3228.740 3377.250 3228.880 ;
        RECT 3368.650 3228.680 3368.970 3228.740 ;
        RECT 3376.930 3228.680 3377.250 3228.740 ;
        RECT 3367.270 3171.760 3367.590 3171.820 ;
        RECT 3369.110 3171.760 3369.430 3171.820 ;
        RECT 3376.930 3171.760 3377.250 3171.820 ;
        RECT 3367.270 3171.620 3377.250 3171.760 ;
        RECT 3367.270 3171.560 3367.590 3171.620 ;
        RECT 3369.110 3171.560 3369.430 3171.620 ;
        RECT 3376.930 3171.560 3377.250 3171.620 ;
      LAYER met1 ;
        RECT 3381.155 3162.855 3588.000 3243.145 ;
      LAYER met1 ;
        RECT 211.210 3118.380 211.530 3118.440 ;
        RECT 213.050 3118.380 213.370 3118.440 ;
        RECT 211.210 3118.240 213.370 3118.380 ;
        RECT 211.210 3118.180 211.530 3118.240 ;
        RECT 213.050 3118.180 213.370 3118.240 ;
        RECT 224.090 3092.000 224.410 3092.260 ;
        RECT 224.180 3091.580 224.320 3092.000 ;
        RECT 224.090 3091.320 224.410 3091.580 ;
        RECT 224.090 3022.500 224.410 3022.560 ;
        RECT 223.720 3022.360 224.410 3022.500 ;
        RECT 223.720 3022.220 223.860 3022.360 ;
        RECT 224.090 3022.300 224.410 3022.360 ;
        RECT 223.630 3021.960 223.950 3022.220 ;
        RECT 221.790 2898.060 222.110 2898.120 ;
        RECT 222.710 2898.060 223.030 2898.120 ;
        RECT 221.790 2897.920 223.030 2898.060 ;
        RECT 221.790 2897.860 222.110 2897.920 ;
        RECT 222.710 2897.860 223.030 2897.920 ;
        RECT 221.790 2801.500 222.110 2801.560 ;
        RECT 223.170 2801.500 223.490 2801.560 ;
        RECT 221.790 2801.360 223.490 2801.500 ;
        RECT 221.790 2801.300 222.110 2801.360 ;
        RECT 223.170 2801.300 223.490 2801.360 ;
      LAYER met1 ;
        RECT 0.000 2557.855 206.845 2638.145 ;
      LAYER met1 ;
        RECT 3369.110 2636.060 3369.430 2636.320 ;
        RECT 3369.200 2635.640 3369.340 2636.060 ;
        RECT 3369.110 2635.380 3369.430 2635.640 ;
        RECT 208.910 2629.460 209.230 2629.520 ;
        RECT 213.050 2629.460 213.370 2629.520 ;
        RECT 208.910 2629.320 213.370 2629.460 ;
        RECT 208.910 2629.260 209.230 2629.320 ;
        RECT 213.050 2629.260 213.370 2629.320 ;
        RECT 3367.270 2614.500 3367.590 2614.560 ;
        RECT 3368.650 2614.500 3368.970 2614.560 ;
        RECT 3376.930 2614.500 3377.250 2614.560 ;
        RECT 3367.270 2614.360 3377.250 2614.500 ;
        RECT 3367.270 2614.300 3367.590 2614.360 ;
        RECT 3368.650 2614.300 3368.970 2614.360 ;
        RECT 3376.930 2614.300 3377.250 2614.360 ;
        RECT 223.630 2608.380 223.950 2608.440 ;
        RECT 224.090 2608.380 224.410 2608.440 ;
        RECT 223.630 2608.240 224.410 2608.380 ;
        RECT 223.630 2608.180 223.950 2608.240 ;
        RECT 224.090 2608.180 224.410 2608.240 ;
        RECT 3369.110 2608.380 3369.430 2608.440 ;
        RECT 3370.030 2608.380 3370.350 2608.440 ;
        RECT 3369.110 2608.240 3370.350 2608.380 ;
        RECT 3369.110 2608.180 3369.430 2608.240 ;
        RECT 3370.030 2608.180 3370.350 2608.240 ;
        RECT 3368.190 2565.540 3368.510 2565.600 ;
        RECT 3370.030 2565.540 3370.350 2565.600 ;
        RECT 3376.930 2565.540 3377.250 2565.600 ;
        RECT 3368.190 2565.400 3377.250 2565.540 ;
        RECT 3368.190 2565.340 3368.510 2565.400 ;
        RECT 3370.030 2565.340 3370.350 2565.400 ;
        RECT 3376.930 2565.340 3377.250 2565.400 ;
      LAYER met1 ;
        RECT 3381.155 2553.855 3588.000 2634.145 ;
      LAYER met1 ;
        RECT 222.710 2521.340 223.030 2521.400 ;
        RECT 223.630 2521.340 223.950 2521.400 ;
        RECT 222.710 2521.200 223.950 2521.340 ;
        RECT 222.710 2521.140 223.030 2521.200 ;
        RECT 223.630 2521.140 223.950 2521.200 ;
        RECT 222.710 2442.460 223.030 2442.520 ;
        RECT 223.630 2442.460 223.950 2442.520 ;
        RECT 222.710 2442.320 223.950 2442.460 ;
        RECT 222.710 2442.260 223.030 2442.320 ;
        RECT 223.630 2442.260 223.950 2442.320 ;
        RECT 223.630 2346.580 223.950 2346.640 ;
        RECT 223.260 2346.440 223.950 2346.580 ;
        RECT 223.260 2345.960 223.400 2346.440 ;
        RECT 223.630 2346.380 223.950 2346.440 ;
        RECT 223.170 2345.700 223.490 2345.960 ;
        RECT 223.170 2318.360 223.490 2318.420 ;
        RECT 224.090 2318.360 224.410 2318.420 ;
        RECT 223.170 2318.220 224.410 2318.360 ;
        RECT 223.170 2318.160 223.490 2318.220 ;
        RECT 224.090 2318.160 224.410 2318.220 ;
        RECT 223.170 2221.800 223.490 2221.860 ;
        RECT 224.090 2221.800 224.410 2221.860 ;
        RECT 223.170 2221.660 224.410 2221.800 ;
        RECT 223.170 2221.600 223.490 2221.660 ;
        RECT 224.090 2221.600 224.410 2221.660 ;
      LAYER met1 ;
        RECT 0.000 1948.855 206.845 2029.145 ;
      LAYER met1 ;
        RECT 208.910 2015.760 209.230 2015.820 ;
        RECT 212.590 2015.760 212.910 2015.820 ;
        RECT 208.910 2015.620 212.910 2015.760 ;
        RECT 208.910 2015.560 209.230 2015.620 ;
        RECT 212.590 2015.560 212.910 2015.620 ;
        RECT 3367.270 2006.920 3367.590 2006.980 ;
        RECT 3369.110 2006.920 3369.430 2006.980 ;
        RECT 3376.930 2006.920 3377.250 2006.980 ;
        RECT 3367.270 2006.780 3377.250 2006.920 ;
        RECT 3367.270 2006.720 3367.590 2006.780 ;
        RECT 3369.110 2006.720 3369.430 2006.780 ;
        RECT 3376.930 2006.720 3377.250 2006.780 ;
        RECT 208.910 1968.500 209.230 1968.560 ;
        RECT 212.130 1968.500 212.450 1968.560 ;
        RECT 208.910 1968.360 212.450 1968.500 ;
        RECT 208.910 1968.300 209.230 1968.360 ;
        RECT 212.130 1968.300 212.450 1968.360 ;
        RECT 224.090 1959.800 224.410 1960.060 ;
        RECT 224.180 1959.380 224.320 1959.800 ;
        RECT 224.090 1959.120 224.410 1959.380 ;
        RECT 3368.190 1958.640 3368.510 1958.700 ;
        RECT 3368.190 1958.500 3377.160 1958.640 ;
        RECT 3368.190 1958.440 3368.510 1958.500 ;
        RECT 3377.020 1958.360 3377.160 1958.500 ;
        RECT 3376.930 1958.100 3377.250 1958.360 ;
      LAYER met1 ;
        RECT 3381.155 1944.855 3588.000 2025.145 ;
      LAYER met1 ;
        RECT 3369.570 1931.780 3369.890 1931.840 ;
        RECT 3370.030 1931.780 3370.350 1931.840 ;
        RECT 3369.570 1931.640 3370.350 1931.780 ;
        RECT 3369.570 1931.580 3369.890 1931.640 ;
        RECT 3370.030 1931.580 3370.350 1931.640 ;
        RECT 223.630 1835.560 223.950 1835.620 ;
        RECT 224.090 1835.560 224.410 1835.620 ;
        RECT 223.630 1835.420 224.410 1835.560 ;
        RECT 223.630 1835.360 223.950 1835.420 ;
        RECT 224.090 1835.360 224.410 1835.420 ;
        RECT 222.250 1738.660 222.570 1738.720 ;
        RECT 224.090 1738.660 224.410 1738.720 ;
        RECT 222.250 1738.520 224.410 1738.660 ;
        RECT 222.250 1738.460 222.570 1738.520 ;
        RECT 224.090 1738.460 224.410 1738.520 ;
        RECT 222.250 1642.440 222.570 1642.500 ;
        RECT 223.630 1642.440 223.950 1642.500 ;
        RECT 222.250 1642.300 223.950 1642.440 ;
        RECT 222.250 1642.240 222.570 1642.300 ;
        RECT 223.630 1642.240 223.950 1642.300 ;
        RECT 222.710 1573.420 223.030 1573.480 ;
        RECT 223.630 1573.420 223.950 1573.480 ;
        RECT 222.710 1573.280 223.950 1573.420 ;
        RECT 222.710 1573.220 223.030 1573.280 ;
        RECT 223.630 1573.220 223.950 1573.280 ;
        RECT 3369.570 1545.880 3369.890 1545.940 ;
        RECT 3370.490 1545.880 3370.810 1545.940 ;
        RECT 3369.570 1545.740 3370.810 1545.880 ;
        RECT 3369.570 1545.680 3369.890 1545.740 ;
        RECT 3370.490 1545.680 3370.810 1545.740 ;
        RECT 222.710 1545.540 223.030 1545.600 ;
        RECT 223.630 1545.540 223.950 1545.600 ;
        RECT 222.710 1545.400 223.950 1545.540 ;
        RECT 222.710 1545.340 223.030 1545.400 ;
        RECT 223.630 1545.340 223.950 1545.400 ;
        RECT 3369.570 1545.200 3369.890 1545.260 ;
        RECT 3370.490 1545.200 3370.810 1545.260 ;
        RECT 3369.570 1545.060 3370.810 1545.200 ;
        RECT 3369.570 1545.000 3369.890 1545.060 ;
        RECT 3370.490 1545.000 3370.810 1545.060 ;
        RECT 222.710 1476.520 223.030 1476.580 ;
        RECT 223.630 1476.520 223.950 1476.580 ;
        RECT 222.710 1476.380 223.950 1476.520 ;
        RECT 222.710 1476.320 223.030 1476.380 ;
        RECT 223.630 1476.320 223.950 1476.380 ;
        RECT 222.710 1448.980 223.030 1449.040 ;
        RECT 224.090 1448.980 224.410 1449.040 ;
        RECT 222.710 1448.840 224.410 1448.980 ;
        RECT 222.710 1448.780 223.030 1448.840 ;
        RECT 224.090 1448.780 224.410 1448.840 ;
      LAYER met1 ;
        RECT 0.000 1340.855 206.845 1421.145 ;
      LAYER met1 ;
        RECT 3369.110 1419.060 3369.430 1419.120 ;
        RECT 3376.470 1419.060 3376.790 1419.120 ;
        RECT 3369.110 1418.920 3376.790 1419.060 ;
        RECT 3369.110 1418.860 3369.430 1418.920 ;
        RECT 3376.470 1418.860 3376.790 1418.920 ;
        RECT 208.910 1407.840 209.230 1407.900 ;
        RECT 212.590 1407.840 212.910 1407.900 ;
        RECT 208.910 1407.700 212.910 1407.840 ;
        RECT 208.910 1407.640 209.230 1407.700 ;
        RECT 212.590 1407.640 212.910 1407.700 ;
        RECT 222.710 1379.620 223.030 1379.680 ;
        RECT 224.090 1379.620 224.410 1379.680 ;
        RECT 222.710 1379.480 224.410 1379.620 ;
        RECT 222.710 1379.420 223.030 1379.480 ;
        RECT 224.090 1379.420 224.410 1379.480 ;
        RECT 208.910 1360.580 209.230 1360.640 ;
        RECT 212.130 1360.580 212.450 1360.640 ;
        RECT 208.910 1360.440 212.450 1360.580 ;
        RECT 208.910 1360.380 209.230 1360.440 ;
        RECT 212.130 1360.380 212.450 1360.440 ;
        RECT 221.790 1352.420 222.110 1352.480 ;
        RECT 222.710 1352.420 223.030 1352.480 ;
        RECT 221.790 1352.280 223.030 1352.420 ;
        RECT 221.790 1352.220 222.110 1352.280 ;
        RECT 222.710 1352.220 223.030 1352.280 ;
        RECT 3369.110 1345.620 3369.430 1345.680 ;
        RECT 3370.490 1345.620 3370.810 1345.680 ;
        RECT 3376.930 1345.620 3377.250 1345.680 ;
        RECT 3369.110 1345.480 3377.250 1345.620 ;
        RECT 3369.110 1345.420 3369.430 1345.480 ;
        RECT 3370.490 1345.420 3370.810 1345.480 ;
        RECT 3376.930 1345.420 3377.250 1345.480 ;
      LAYER met1 ;
        RECT 3381.155 1336.855 3588.000 1417.145 ;
      LAYER met1 ;
        RECT 221.790 1256.200 222.110 1256.260 ;
        RECT 223.170 1256.200 223.490 1256.260 ;
        RECT 221.790 1256.060 223.490 1256.200 ;
        RECT 221.790 1256.000 222.110 1256.060 ;
        RECT 223.170 1256.000 223.490 1256.060 ;
        RECT 223.630 1062.740 223.950 1062.800 ;
        RECT 224.090 1062.740 224.410 1062.800 ;
        RECT 223.630 1062.600 224.410 1062.740 ;
        RECT 223.630 1062.540 223.950 1062.600 ;
        RECT 224.090 1062.540 224.410 1062.600 ;
        RECT 223.630 897.160 223.950 897.220 ;
        RECT 223.260 897.020 223.950 897.160 ;
        RECT 223.260 896.880 223.400 897.020 ;
        RECT 223.630 896.960 223.950 897.020 ;
        RECT 3368.650 897.160 3368.970 897.220 ;
        RECT 3369.570 897.160 3369.890 897.220 ;
        RECT 3368.650 897.020 3369.890 897.160 ;
        RECT 3368.650 896.960 3368.970 897.020 ;
        RECT 3369.570 896.960 3369.890 897.020 ;
        RECT 223.170 896.620 223.490 896.880 ;
        RECT 223.170 869.620 223.490 869.680 ;
        RECT 223.630 869.620 223.950 869.680 ;
        RECT 223.170 869.480 223.950 869.620 ;
        RECT 223.170 869.420 223.490 869.480 ;
        RECT 223.630 869.420 223.950 869.480 ;
      LAYER met1 ;
        RECT 0.000 731.855 206.845 812.145 ;
      LAYER met1 ;
        RECT 208.910 800.260 209.230 800.320 ;
        RECT 212.590 800.260 212.910 800.320 ;
        RECT 208.910 800.120 212.910 800.260 ;
        RECT 208.910 800.060 209.230 800.120 ;
        RECT 212.590 800.060 212.910 800.120 ;
        RECT 3368.190 788.700 3368.510 788.760 ;
        RECT 3376.930 788.700 3377.250 788.760 ;
        RECT 3368.190 788.560 3377.250 788.700 ;
        RECT 3368.190 788.500 3368.510 788.560 ;
        RECT 3376.930 788.500 3377.250 788.560 ;
        RECT 208.910 750.960 209.230 751.020 ;
        RECT 212.130 750.960 212.450 751.020 ;
        RECT 208.910 750.820 212.450 750.960 ;
        RECT 208.910 750.760 209.230 750.820 ;
        RECT 212.130 750.760 212.450 750.820 ;
        RECT 3367.270 741.440 3367.590 741.500 ;
        RECT 3368.650 741.440 3368.970 741.500 ;
        RECT 3376.930 741.440 3377.250 741.500 ;
        RECT 3367.270 741.300 3377.250 741.440 ;
        RECT 3367.270 741.240 3367.590 741.300 ;
        RECT 3368.650 741.240 3368.970 741.300 ;
        RECT 3376.930 741.240 3377.250 741.300 ;
      LAYER met1 ;
        RECT 3381.155 727.855 3588.000 808.145 ;
      LAYER met1 ;
        RECT 223.170 579.940 223.490 580.000 ;
        RECT 223.170 579.800 223.860 579.940 ;
        RECT 223.170 579.740 223.490 579.800 ;
        RECT 223.720 578.980 223.860 579.800 ;
        RECT 223.630 578.720 223.950 578.980 ;
        RECT 224.090 386.960 224.410 387.220 ;
        RECT 224.180 386.540 224.320 386.960 ;
        RECT 224.090 386.280 224.410 386.540 ;
        RECT 2911.870 228.720 2912.190 228.780 ;
        RECT 3373.710 228.720 3374.030 228.780 ;
        RECT 2911.870 228.580 3374.030 228.720 ;
        RECT 2911.870 228.520 2912.190 228.580 ;
        RECT 3373.710 228.520 3374.030 228.580 ;
        RECT 212.130 228.380 212.450 228.440 ;
        RECT 1257.710 228.380 1258.030 228.440 ;
        RECT 212.130 228.240 1258.030 228.380 ;
        RECT 212.130 228.180 212.450 228.240 ;
        RECT 1257.710 228.180 1258.030 228.240 ;
        RECT 2348.830 228.380 2349.150 228.440 ;
        RECT 3367.270 228.380 3367.590 228.440 ;
        RECT 2348.830 228.240 3367.590 228.380 ;
        RECT 2348.830 228.180 2349.150 228.240 ;
        RECT 3367.270 228.180 3367.590 228.240 ;
        RECT 2370.450 228.040 2370.770 228.100 ;
        RECT 3368.190 228.040 3368.510 228.100 ;
        RECT 2370.450 227.900 3368.510 228.040 ;
        RECT 2370.450 227.840 2370.770 227.900 ;
        RECT 3368.190 227.840 3368.510 227.900 ;
        RECT 224.550 227.700 224.870 227.760 ;
        RECT 1800.050 227.700 1800.370 227.760 ;
        RECT 224.550 227.560 1800.370 227.700 ;
        RECT 224.550 227.500 224.870 227.560 ;
        RECT 1800.050 227.500 1800.370 227.560 ;
        RECT 741.130 221.920 741.450 221.980 ;
        RECT 1815.230 221.920 1815.550 221.980 ;
        RECT 1821.210 221.920 1821.530 221.980 ;
        RECT 741.130 221.780 1821.530 221.920 ;
        RECT 741.130 221.720 741.450 221.780 ;
        RECT 1815.230 221.720 1815.550 221.780 ;
        RECT 1821.210 221.720 1821.530 221.780 ;
        RECT 1824.430 221.920 1824.750 221.980 ;
        RECT 2304.670 221.920 2304.990 221.980 ;
        RECT 1824.430 221.780 2304.990 221.920 ;
        RECT 1824.430 221.720 1824.750 221.780 ;
        RECT 2304.670 221.720 2304.990 221.780 ;
        RECT 1827.650 221.580 1827.970 221.640 ;
        RECT 2325.370 221.580 2325.690 221.640 ;
        RECT 2348.830 221.580 2349.150 221.640 ;
        RECT 1827.650 221.440 2349.150 221.580 ;
        RECT 1827.650 221.380 1827.970 221.440 ;
        RECT 2325.370 221.380 2325.690 221.440 ;
        RECT 2348.830 221.380 2349.150 221.440 ;
        RECT 1257.710 221.240 1258.030 221.300 ;
        RECT 2353.430 221.240 2353.750 221.300 ;
        RECT 2370.450 221.240 2370.770 221.300 ;
        RECT 1257.710 221.100 2370.770 221.240 ;
        RECT 1257.710 221.040 1258.030 221.100 ;
        RECT 2353.430 221.040 2353.750 221.100 ;
        RECT 2370.450 221.040 2370.770 221.100 ;
        RECT 1821.210 220.900 1821.530 220.960 ;
        RECT 2332.270 220.900 2332.590 220.960 ;
        RECT 2891.630 220.900 2891.950 220.960 ;
        RECT 2911.870 220.900 2912.190 220.960 ;
        RECT 1821.210 220.760 2912.190 220.900 ;
        RECT 1821.210 220.700 1821.530 220.760 ;
        RECT 2332.270 220.700 2332.590 220.760 ;
        RECT 2891.630 220.700 2891.950 220.760 ;
        RECT 2911.870 220.700 2912.190 220.760 ;
        RECT 212.590 213.760 212.910 213.820 ;
        RECT 1283.010 213.760 1283.330 213.820 ;
        RECT 212.590 213.620 1283.330 213.760 ;
        RECT 212.590 213.560 212.910 213.620 ;
        RECT 1283.010 213.560 1283.330 213.620 ;
        RECT 1784.870 211.380 1785.190 211.440 ;
        RECT 1827.650 211.380 1827.970 211.440 ;
        RECT 1784.870 211.240 1827.970 211.380 ;
        RECT 1784.870 211.180 1785.190 211.240 ;
        RECT 1827.650 211.180 1827.970 211.240 ;
        RECT 1784.870 209.340 1785.190 209.400 ;
        RECT 1763.340 209.200 1785.190 209.340 ;
        RECT 1763.340 209.060 1763.480 209.200 ;
        RECT 1784.870 209.140 1785.190 209.200 ;
        RECT 1812.470 209.340 1812.790 209.400 ;
        RECT 1820.290 209.340 1820.610 209.400 ;
        RECT 1812.470 209.200 1820.610 209.340 ;
        RECT 1812.470 209.140 1812.790 209.200 ;
        RECT 1820.290 209.140 1820.610 209.200 ;
        RECT 1763.250 208.800 1763.570 209.060 ;
        RECT 1766.470 209.000 1766.790 209.060 ;
        RECT 1774.290 209.000 1774.610 209.060 ;
        RECT 1780.270 209.000 1780.590 209.060 ;
        RECT 1786.710 209.000 1787.030 209.060 ;
        RECT 1801.890 209.000 1802.210 209.060 ;
        RECT 1766.470 208.860 1802.210 209.000 ;
        RECT 1766.470 208.800 1766.790 208.860 ;
        RECT 1774.290 208.800 1774.610 208.860 ;
        RECT 1780.270 208.800 1780.590 208.860 ;
        RECT 1786.710 208.800 1787.030 208.860 ;
        RECT 1801.890 208.800 1802.210 208.860 ;
        RECT 1283.010 207.640 1283.330 207.700 ;
        RECT 1379.610 207.640 1379.930 207.700 ;
        RECT 1283.010 207.500 1379.930 207.640 ;
        RECT 1283.010 207.440 1283.330 207.500 ;
        RECT 1379.610 207.440 1379.930 207.500 ;
        RECT 1380.070 207.640 1380.390 207.700 ;
        RECT 1545.210 207.640 1545.530 207.700 ;
        RECT 1572.810 207.640 1573.130 207.700 ;
        RECT 1380.070 207.500 1400.540 207.640 ;
        RECT 1380.070 207.440 1380.390 207.500 ;
        RECT 1400.400 207.300 1400.540 207.500 ;
        RECT 1545.210 207.500 1573.130 207.640 ;
        RECT 1545.210 207.440 1545.530 207.500 ;
        RECT 1572.810 207.440 1573.130 207.500 ;
        RECT 1573.270 207.640 1573.590 207.700 ;
        RECT 1573.270 207.500 1593.740 207.640 ;
        RECT 1573.270 207.440 1573.590 207.500 ;
        RECT 1449.070 207.300 1449.390 207.360 ;
        RECT 1400.400 207.160 1449.390 207.300 ;
        RECT 1593.600 207.300 1593.740 207.500 ;
        RECT 1642.270 207.300 1642.590 207.360 ;
        RECT 1593.600 207.160 1642.590 207.300 ;
        RECT 1449.070 207.100 1449.390 207.160 ;
        RECT 1642.270 207.100 1642.590 207.160 ;
        RECT 1711.270 207.300 1711.590 207.360 ;
        RECT 1763.340 207.300 1763.480 208.800 ;
        RECT 1711.270 207.160 1763.480 207.300 ;
        RECT 1711.270 207.100 1711.590 207.160 ;
        RECT 1211.480 200.840 1211.800 200.900 ;
        RECT 1265.070 200.840 1265.390 200.900 ;
        RECT 1211.480 200.700 1265.390 200.840 ;
        RECT 1211.480 200.640 1211.800 200.700 ;
        RECT 1265.070 200.640 1265.390 200.700 ;
        RECT 1257.710 200.500 1258.030 200.560 ;
        RECT 1262.770 200.500 1263.090 200.560 ;
        RECT 1250.900 200.360 1268.980 200.500 ;
        RECT 1250.900 200.000 1251.040 200.360 ;
        RECT 1257.710 200.300 1258.030 200.360 ;
        RECT 1258.950 200.000 1259.090 200.360 ;
        RECT 1261.430 200.000 1261.570 200.360 ;
        RECT 1262.770 200.300 1263.090 200.360 ;
        RECT 1268.840 200.000 1268.980 200.360 ;
      LAYER met1 ;
        RECT 668.380 0.275 741.815 197.965 ;
        RECT 1209.000 189.745 1258.585 200.000 ;
      LAYER met1 ;
        RECT 1258.865 190.025 1259.095 200.000 ;
      LAYER met1 ;
        RECT 1259.375 189.745 1284.000 200.000 ;
        RECT 1209.000 0.790 1284.000 189.745 ;
        RECT 1751.855 0.000 1832.145 206.845 ;
      LAYER met1 ;
        RECT 2299.150 198.460 2299.470 198.520 ;
        RECT 2304.670 198.460 2304.990 198.520 ;
        RECT 2299.150 198.320 2304.990 198.460 ;
        RECT 2299.150 198.260 2299.470 198.320 ;
        RECT 2304.670 198.260 2304.990 198.320 ;
      LAYER met1 ;
        RECT 2299.215 0.160 2373.880 197.965 ;
        RECT 2843.085 0.275 2915.815 197.965 ;
      LAYER via ;
        RECT 707.120 4977.980 707.380 4978.240 ;
        RECT 745.760 4977.980 746.020 4978.240 ;
        RECT 2341.960 4977.300 2342.220 4977.560 ;
        RECT 2380.600 4977.300 2380.860 4977.560 ;
        RECT 1251.760 4976.960 1252.020 4977.220 ;
        RECT 1290.860 4976.960 1291.120 4977.220 ;
        RECT 1228.300 4960.300 1228.560 4960.560 ;
        RECT 1282.120 4960.300 1282.380 4960.560 ;
        RECT 684.580 4953.840 684.840 4954.100 ;
        RECT 1226.000 4953.840 1226.260 4954.100 ;
        RECT 1796.400 4953.840 1796.660 4954.100 ;
        RECT 1836.420 4953.840 1836.680 4954.100 ;
        RECT 1827.220 4953.500 1827.480 4953.760 ;
        RECT 2370.020 4953.840 2370.280 4954.100 ;
        RECT 2372.320 4953.840 2372.580 4954.100 ;
        RECT 1089.840 4953.160 1090.100 4953.420 ;
        RECT 224.120 4952.140 224.380 4952.400 ;
        RECT 317.500 4952.140 317.760 4952.400 ;
        RECT 412.260 4952.140 412.520 4952.400 ;
        RECT 662.500 4952.480 662.760 4952.740 ;
        RECT 737.020 4952.480 737.280 4952.740 ;
        RECT 1282.120 4952.480 1282.380 4952.740 ;
        RECT 1435.300 4952.480 1435.560 4952.740 ;
        RECT 1545.240 4952.480 1545.500 4952.740 ;
        RECT 1628.500 4952.480 1628.760 4952.740 ;
        RECT 1738.440 4952.480 1738.700 4952.740 ;
        RECT 1827.220 4952.480 1827.480 4952.740 ;
        RECT 224.580 4951.460 224.840 4951.720 ;
        RECT 386.500 4951.120 386.760 4951.380 ;
        RECT 530.940 4951.800 531.200 4952.060 ;
        RECT 772.900 4952.140 773.160 4952.400 ;
        RECT 1226.000 4952.140 1226.260 4952.400 ;
        RECT 1229.680 4952.140 1229.940 4952.400 ;
        RECT 1448.640 4952.140 1448.900 4952.400 ;
        RECT 1449.560 4952.140 1449.820 4952.400 ;
        RECT 1774.780 4952.140 1775.040 4952.400 ;
        RECT 2319.880 4953.500 2320.140 4953.760 ;
        RECT 2856.700 4953.500 2856.960 4953.760 ;
        RECT 758.640 4951.800 758.900 4952.060 ;
        RECT 1179.540 4951.800 1179.800 4952.060 ;
        RECT 1227.840 4951.800 1228.100 4952.060 ;
        RECT 1450.020 4951.800 1450.280 4952.060 ;
        RECT 1545.240 4951.800 1545.500 4952.060 ;
        RECT 317.500 4950.780 317.760 4951.040 ;
        RECT 412.260 4950.780 412.520 4951.040 ;
        RECT 211.240 4950.440 211.500 4950.700 ;
        RECT 414.100 4950.440 414.360 4950.700 ;
        RECT 662.960 4951.120 663.220 4951.380 ;
        RECT 758.640 4951.120 758.900 4951.380 ;
        RECT 684.580 4950.780 684.840 4951.040 ;
        RECT 773.360 4950.780 773.620 4951.040 ;
        RECT 510.700 4950.440 510.960 4950.700 ;
        RECT 530.940 4950.440 531.200 4950.700 ;
        RECT 531.400 4950.440 531.660 4950.700 ;
        RECT 737.020 4950.440 737.280 4950.700 ;
        RECT 966.100 4951.120 966.360 4951.380 ;
        RECT 1089.840 4951.120 1090.100 4951.380 ;
        RECT 1227.380 4951.120 1227.640 4951.380 ;
        RECT 1228.300 4951.120 1228.560 4951.380 ;
        RECT 1380.100 4951.120 1380.360 4951.380 ;
        RECT 1474.860 4951.120 1475.120 4951.380 ;
        RECT 1226.920 4950.780 1227.180 4951.040 ;
        RECT 1227.840 4950.780 1228.100 4951.040 ;
        RECT 1379.640 4950.780 1379.900 4951.040 ;
        RECT 2856.700 4950.780 2856.960 4951.040 ;
        RECT 2870.040 4950.780 2870.300 4951.040 ;
        RECT 3373.740 4950.780 3374.000 4951.040 ;
        RECT 1091.220 4950.440 1091.480 4950.700 ;
        RECT 1179.540 4950.440 1179.800 4950.700 ;
        RECT 2370.020 4950.440 2370.280 4950.700 ;
        RECT 3365.460 4950.440 3365.720 4950.700 ;
        RECT 222.280 4574.400 222.540 4574.660 ;
        RECT 224.120 4574.400 224.380 4574.660 ;
        RECT 3368.680 4471.380 3368.940 4471.640 ;
        RECT 3373.740 4471.380 3374.000 4471.640 ;
        RECT 3390.300 4471.380 3390.560 4471.640 ;
        RECT 222.280 4443.500 222.540 4443.760 ;
        RECT 223.660 4443.500 223.920 4443.760 ;
        RECT 3365.460 4399.980 3365.720 4400.240 ;
        RECT 3368.220 4399.980 3368.480 4400.240 ;
        RECT 3368.220 4380.600 3368.480 4380.860 ;
        RECT 3389.380 4380.600 3389.640 4380.860 ;
        RECT 3373.740 4374.480 3374.000 4374.740 ;
        RECT 3388.460 4374.480 3388.720 4374.740 ;
        RECT 210.780 4346.940 211.040 4347.200 ;
        RECT 223.660 4346.940 223.920 4347.200 ;
        RECT 223.660 4181.360 223.920 4181.620 ;
        RECT 223.200 4181.020 223.460 4181.280 ;
        RECT 223.200 4153.820 223.460 4154.080 ;
        RECT 223.660 4153.820 223.920 4154.080 ;
        RECT 222.280 3891.680 222.540 3891.940 ;
        RECT 222.740 3891.000 223.000 3891.260 ;
        RECT 211.240 3871.280 211.500 3871.540 ;
        RECT 212.620 3871.280 212.880 3871.540 ;
        RECT 208.940 3846.120 209.200 3846.380 ;
        RECT 212.620 3846.120 212.880 3846.380 ;
        RECT 211.700 3836.600 211.960 3836.860 ;
        RECT 212.620 3836.600 212.880 3836.860 ;
        RECT 3368.680 3836.600 3368.940 3836.860 ;
        RECT 3376.960 3836.600 3377.220 3836.860 ;
        RECT 208.940 3792.400 209.200 3792.660 ;
        RECT 213.080 3792.400 213.340 3792.660 ;
        RECT 220.900 3792.400 221.160 3792.660 ;
        RECT 3367.300 3779.480 3367.560 3779.740 ;
        RECT 3368.220 3779.480 3368.480 3779.740 ;
        RECT 3376.960 3779.480 3377.220 3779.740 ;
        RECT 211.700 3757.720 211.960 3757.980 ;
        RECT 213.080 3757.720 213.340 3757.980 ;
        RECT 223.660 3698.560 223.920 3698.820 ;
        RECT 224.120 3697.880 224.380 3698.140 ;
        RECT 223.200 3670.340 223.460 3670.600 ;
        RECT 224.120 3670.340 224.380 3670.600 ;
        RECT 223.200 3601.660 223.460 3601.920 ;
        RECT 224.120 3601.660 224.380 3601.920 ;
        RECT 224.120 3505.100 224.380 3505.360 ;
        RECT 224.120 3504.420 224.380 3504.680 ;
        RECT 222.280 3463.620 222.540 3463.880 ;
        RECT 224.120 3463.620 224.380 3463.880 ;
        RECT 222.280 3367.400 222.540 3367.660 ;
        RECT 223.660 3367.400 223.920 3367.660 ;
        RECT 223.660 3312.320 223.920 3312.580 ;
        RECT 223.200 3311.640 223.460 3311.900 ;
        RECT 211.240 3254.520 211.500 3254.780 ;
        RECT 212.160 3254.520 212.420 3254.780 ;
        RECT 208.940 3238.200 209.200 3238.460 ;
        RECT 212.160 3238.200 212.420 3238.460 ;
        RECT 213.080 3238.200 213.340 3238.460 ;
        RECT 3368.680 3228.680 3368.940 3228.940 ;
        RECT 3376.960 3228.680 3377.220 3228.940 ;
        RECT 3367.300 3171.560 3367.560 3171.820 ;
        RECT 3369.140 3171.560 3369.400 3171.820 ;
        RECT 3376.960 3171.560 3377.220 3171.820 ;
        RECT 211.240 3118.180 211.500 3118.440 ;
        RECT 213.080 3118.180 213.340 3118.440 ;
        RECT 224.120 3092.000 224.380 3092.260 ;
        RECT 224.120 3091.320 224.380 3091.580 ;
        RECT 224.120 3022.300 224.380 3022.560 ;
        RECT 223.660 3021.960 223.920 3022.220 ;
        RECT 221.820 2897.860 222.080 2898.120 ;
        RECT 222.740 2897.860 223.000 2898.120 ;
        RECT 221.820 2801.300 222.080 2801.560 ;
        RECT 223.200 2801.300 223.460 2801.560 ;
        RECT 3369.140 2636.060 3369.400 2636.320 ;
        RECT 3369.140 2635.380 3369.400 2635.640 ;
        RECT 208.940 2629.260 209.200 2629.520 ;
        RECT 213.080 2629.260 213.340 2629.520 ;
        RECT 3367.300 2614.300 3367.560 2614.560 ;
        RECT 3368.680 2614.300 3368.940 2614.560 ;
        RECT 3376.960 2614.300 3377.220 2614.560 ;
        RECT 223.660 2608.180 223.920 2608.440 ;
        RECT 224.120 2608.180 224.380 2608.440 ;
        RECT 3369.140 2608.180 3369.400 2608.440 ;
        RECT 3370.060 2608.180 3370.320 2608.440 ;
        RECT 3368.220 2565.340 3368.480 2565.600 ;
        RECT 3370.060 2565.340 3370.320 2565.600 ;
        RECT 3376.960 2565.340 3377.220 2565.600 ;
        RECT 222.740 2521.140 223.000 2521.400 ;
        RECT 223.660 2521.140 223.920 2521.400 ;
        RECT 222.740 2442.260 223.000 2442.520 ;
        RECT 223.660 2442.260 223.920 2442.520 ;
        RECT 223.660 2346.380 223.920 2346.640 ;
        RECT 223.200 2345.700 223.460 2345.960 ;
        RECT 223.200 2318.160 223.460 2318.420 ;
        RECT 224.120 2318.160 224.380 2318.420 ;
        RECT 223.200 2221.600 223.460 2221.860 ;
        RECT 224.120 2221.600 224.380 2221.860 ;
        RECT 208.940 2015.560 209.200 2015.820 ;
        RECT 212.620 2015.560 212.880 2015.820 ;
        RECT 3367.300 2006.720 3367.560 2006.980 ;
        RECT 3369.140 2006.720 3369.400 2006.980 ;
        RECT 3376.960 2006.720 3377.220 2006.980 ;
        RECT 208.940 1968.300 209.200 1968.560 ;
        RECT 212.160 1968.300 212.420 1968.560 ;
        RECT 224.120 1959.800 224.380 1960.060 ;
        RECT 224.120 1959.120 224.380 1959.380 ;
        RECT 3368.220 1958.440 3368.480 1958.700 ;
        RECT 3376.960 1958.100 3377.220 1958.360 ;
        RECT 3369.600 1931.580 3369.860 1931.840 ;
        RECT 3370.060 1931.580 3370.320 1931.840 ;
        RECT 223.660 1835.360 223.920 1835.620 ;
        RECT 224.120 1835.360 224.380 1835.620 ;
        RECT 222.280 1738.460 222.540 1738.720 ;
        RECT 224.120 1738.460 224.380 1738.720 ;
        RECT 222.280 1642.240 222.540 1642.500 ;
        RECT 223.660 1642.240 223.920 1642.500 ;
        RECT 222.740 1573.220 223.000 1573.480 ;
        RECT 223.660 1573.220 223.920 1573.480 ;
        RECT 3369.600 1545.680 3369.860 1545.940 ;
        RECT 3370.520 1545.680 3370.780 1545.940 ;
        RECT 222.740 1545.340 223.000 1545.600 ;
        RECT 223.660 1545.340 223.920 1545.600 ;
        RECT 3369.600 1545.000 3369.860 1545.260 ;
        RECT 3370.520 1545.000 3370.780 1545.260 ;
        RECT 222.740 1476.320 223.000 1476.580 ;
        RECT 223.660 1476.320 223.920 1476.580 ;
        RECT 222.740 1448.780 223.000 1449.040 ;
        RECT 224.120 1448.780 224.380 1449.040 ;
        RECT 3369.140 1418.860 3369.400 1419.120 ;
        RECT 3376.500 1418.860 3376.760 1419.120 ;
        RECT 208.940 1407.640 209.200 1407.900 ;
        RECT 212.620 1407.640 212.880 1407.900 ;
        RECT 222.740 1379.420 223.000 1379.680 ;
        RECT 224.120 1379.420 224.380 1379.680 ;
        RECT 208.940 1360.380 209.200 1360.640 ;
        RECT 212.160 1360.380 212.420 1360.640 ;
        RECT 221.820 1352.220 222.080 1352.480 ;
        RECT 222.740 1352.220 223.000 1352.480 ;
        RECT 3369.140 1345.420 3369.400 1345.680 ;
        RECT 3370.520 1345.420 3370.780 1345.680 ;
        RECT 3376.960 1345.420 3377.220 1345.680 ;
        RECT 221.820 1256.000 222.080 1256.260 ;
        RECT 223.200 1256.000 223.460 1256.260 ;
        RECT 223.660 1062.540 223.920 1062.800 ;
        RECT 224.120 1062.540 224.380 1062.800 ;
        RECT 223.660 896.960 223.920 897.220 ;
        RECT 3368.680 896.960 3368.940 897.220 ;
        RECT 3369.600 896.960 3369.860 897.220 ;
        RECT 223.200 896.620 223.460 896.880 ;
        RECT 223.200 869.420 223.460 869.680 ;
        RECT 223.660 869.420 223.920 869.680 ;
        RECT 208.940 800.060 209.200 800.320 ;
        RECT 212.620 800.060 212.880 800.320 ;
        RECT 3368.220 788.500 3368.480 788.760 ;
        RECT 3376.960 788.500 3377.220 788.760 ;
        RECT 208.940 750.760 209.200 751.020 ;
        RECT 212.160 750.760 212.420 751.020 ;
        RECT 3367.300 741.240 3367.560 741.500 ;
        RECT 3368.680 741.240 3368.940 741.500 ;
        RECT 3376.960 741.240 3377.220 741.500 ;
        RECT 223.200 579.740 223.460 580.000 ;
        RECT 223.660 578.720 223.920 578.980 ;
        RECT 224.120 386.960 224.380 387.220 ;
        RECT 224.120 386.280 224.380 386.540 ;
        RECT 2911.900 228.520 2912.160 228.780 ;
        RECT 3373.740 228.520 3374.000 228.780 ;
        RECT 212.160 228.180 212.420 228.440 ;
        RECT 1257.740 228.180 1258.000 228.440 ;
        RECT 2348.860 228.180 2349.120 228.440 ;
        RECT 3367.300 228.180 3367.560 228.440 ;
        RECT 2370.480 227.840 2370.740 228.100 ;
        RECT 3368.220 227.840 3368.480 228.100 ;
        RECT 224.580 227.500 224.840 227.760 ;
        RECT 1800.080 227.500 1800.340 227.760 ;
        RECT 741.160 221.720 741.420 221.980 ;
        RECT 1815.260 221.720 1815.520 221.980 ;
        RECT 1821.240 221.720 1821.500 221.980 ;
        RECT 1824.460 221.720 1824.720 221.980 ;
        RECT 2304.700 221.720 2304.960 221.980 ;
        RECT 1827.680 221.380 1827.940 221.640 ;
        RECT 2325.400 221.380 2325.660 221.640 ;
        RECT 2348.860 221.380 2349.120 221.640 ;
        RECT 1257.740 221.040 1258.000 221.300 ;
        RECT 2353.460 221.040 2353.720 221.300 ;
        RECT 2370.480 221.040 2370.740 221.300 ;
        RECT 1821.240 220.700 1821.500 220.960 ;
        RECT 2332.300 220.700 2332.560 220.960 ;
        RECT 2891.660 220.700 2891.920 220.960 ;
        RECT 2911.900 220.700 2912.160 220.960 ;
        RECT 212.620 213.560 212.880 213.820 ;
        RECT 1283.040 213.560 1283.300 213.820 ;
        RECT 1784.900 211.180 1785.160 211.440 ;
        RECT 1827.680 211.180 1827.940 211.440 ;
        RECT 1784.900 209.140 1785.160 209.400 ;
        RECT 1812.500 209.140 1812.760 209.400 ;
        RECT 1820.320 209.140 1820.580 209.400 ;
        RECT 1763.280 208.800 1763.540 209.060 ;
        RECT 1766.500 208.800 1766.760 209.060 ;
        RECT 1774.320 208.800 1774.580 209.060 ;
        RECT 1780.300 208.800 1780.560 209.060 ;
        RECT 1786.740 208.800 1787.000 209.060 ;
        RECT 1801.920 208.800 1802.180 209.060 ;
        RECT 1283.040 207.440 1283.300 207.700 ;
        RECT 1379.640 207.440 1379.900 207.700 ;
        RECT 1380.100 207.440 1380.360 207.700 ;
        RECT 1545.240 207.440 1545.500 207.700 ;
        RECT 1572.840 207.440 1573.100 207.700 ;
        RECT 1573.300 207.440 1573.560 207.700 ;
        RECT 1449.100 207.100 1449.360 207.360 ;
        RECT 1642.300 207.100 1642.560 207.360 ;
        RECT 1711.300 207.100 1711.560 207.360 ;
        RECT 1211.510 200.640 1211.770 200.900 ;
        RECT 1265.100 200.640 1265.360 200.900 ;
        RECT 1257.740 200.300 1258.000 200.560 ;
        RECT 1262.800 200.300 1263.060 200.560 ;
        RECT 2299.180 198.260 2299.440 198.520 ;
        RECT 2304.700 198.260 2304.960 198.520 ;
      LAYER met2 ;
        RECT 668.210 4979.715 747.915 5188.000 ;
        RECT 668.210 4979.435 669.205 4979.715 ;
        RECT 670.045 4979.435 671.965 4979.715 ;
        RECT 672.805 4979.435 675.185 4979.715 ;
        RECT 676.025 4979.435 678.405 4979.715 ;
        RECT 679.245 4979.435 681.165 4979.715 ;
        RECT 682.005 4979.435 684.385 4979.715 ;
        RECT 685.225 4979.435 687.605 4979.715 ;
        RECT 688.445 4979.435 690.365 4979.715 ;
        RECT 691.205 4979.435 693.585 4979.715 ;
        RECT 694.425 4979.435 696.805 4979.715 ;
        RECT 697.645 4979.435 699.565 4979.715 ;
        RECT 700.405 4979.435 702.785 4979.715 ;
        RECT 703.625 4979.435 706.005 4979.715 ;
        RECT 706.845 4979.435 709.225 4979.715 ;
        RECT 710.065 4979.435 711.985 4979.715 ;
        RECT 712.825 4979.435 715.205 4979.715 ;
        RECT 716.045 4979.435 718.425 4979.715 ;
        RECT 719.265 4979.435 721.185 4979.715 ;
        RECT 722.025 4979.435 724.405 4979.715 ;
        RECT 725.245 4979.435 727.625 4979.715 ;
        RECT 728.465 4979.435 730.385 4979.715 ;
        RECT 731.225 4979.435 733.605 4979.715 ;
        RECT 734.445 4979.435 736.825 4979.715 ;
        RECT 737.665 4979.435 739.585 4979.715 ;
        RECT 740.425 4979.435 742.805 4979.715 ;
        RECT 743.645 4979.435 746.025 4979.715 ;
        RECT 746.865 4979.435 747.915 4979.715 ;
        RECT 1213.210 4979.715 1292.915 5188.000 ;
      LAYER met2 ;
        RECT 1620.210 4982.515 1620.490 4982.885 ;
      LAYER met2 ;
        RECT 1213.210 4979.435 1214.205 4979.715 ;
        RECT 1215.045 4979.435 1216.965 4979.715 ;
        RECT 1217.805 4979.435 1220.185 4979.715 ;
        RECT 1221.025 4979.435 1223.405 4979.715 ;
        RECT 1224.245 4979.435 1226.165 4979.715 ;
        RECT 1227.005 4979.435 1229.385 4979.715 ;
        RECT 1230.225 4979.435 1232.605 4979.715 ;
        RECT 1233.445 4979.435 1235.365 4979.715 ;
        RECT 1236.205 4979.435 1238.585 4979.715 ;
        RECT 1239.425 4979.435 1241.805 4979.715 ;
        RECT 1242.645 4979.435 1244.565 4979.715 ;
        RECT 1245.405 4979.435 1247.785 4979.715 ;
        RECT 1248.625 4979.435 1251.005 4979.715 ;
        RECT 1251.845 4979.435 1254.225 4979.715 ;
        RECT 1255.065 4979.435 1256.985 4979.715 ;
        RECT 1257.825 4979.435 1260.205 4979.715 ;
        RECT 1261.045 4979.435 1263.425 4979.715 ;
        RECT 1264.265 4979.435 1266.185 4979.715 ;
        RECT 1267.025 4979.435 1269.405 4979.715 ;
        RECT 1270.245 4979.435 1272.625 4979.715 ;
        RECT 1273.465 4979.435 1275.385 4979.715 ;
        RECT 1276.225 4979.435 1278.605 4979.715 ;
        RECT 1279.445 4979.435 1281.825 4979.715 ;
        RECT 1282.665 4979.435 1284.585 4979.715 ;
        RECT 1285.425 4979.435 1287.805 4979.715 ;
        RECT 1288.645 4979.435 1291.025 4979.715 ;
        RECT 1291.865 4979.435 1292.915 4979.715 ;
      LAYER met2 ;
        RECT 669.485 4977.035 669.765 4979.435 ;
        RECT 684.665 4977.260 684.945 4979.435 ;
        RECT 684.640 4977.035 684.945 4977.260 ;
        RECT 706.285 4977.330 706.565 4979.435 ;
        RECT 707.120 4977.950 707.380 4978.270 ;
        RECT 707.180 4977.330 707.320 4977.950 ;
        RECT 706.285 4977.190 707.320 4977.330 ;
        RECT 706.285 4977.035 706.565 4977.190 ;
        RECT 721.465 4977.035 721.745 4979.435 ;
        RECT 727.905 4977.035 728.185 4979.435 ;
        RECT 730.665 4977.035 730.945 4979.435 ;
        RECT 737.105 4977.260 737.385 4979.435 ;
        RECT 737.080 4977.035 737.385 4977.260 ;
        RECT 739.865 4977.035 740.145 4979.435 ;
        RECT 746.305 4978.305 746.585 4979.435 ;
        RECT 745.820 4978.270 746.585 4978.305 ;
        RECT 745.760 4978.165 746.585 4978.270 ;
        RECT 745.760 4977.950 746.020 4978.165 ;
        RECT 746.305 4977.035 746.585 4978.165 ;
        RECT 1214.485 4977.035 1214.765 4979.435 ;
        RECT 1229.665 4977.035 1229.945 4979.435 ;
        RECT 1251.285 4977.330 1251.565 4979.435 ;
        RECT 1251.285 4977.250 1251.960 4977.330 ;
        RECT 1251.285 4977.190 1252.020 4977.250 ;
        RECT 1251.285 4977.035 1251.565 4977.190 ;
        RECT 684.640 4954.130 684.780 4977.035 ;
        RECT 684.580 4953.810 684.840 4954.130 ;
        RECT 662.560 4952.770 663.160 4952.850 ;
        RECT 662.500 4952.710 663.160 4952.770 ;
        RECT 662.500 4952.450 662.760 4952.710 ;
        RECT 224.120 4952.110 224.380 4952.430 ;
        RECT 317.500 4952.110 317.760 4952.430 ;
        RECT 412.260 4952.110 412.520 4952.430 ;
        RECT 211.240 4950.410 211.500 4950.730 ;
      LAYER met2 ;
        RECT 4.925 4434.110 174.060 4458.290 ;
      LAYER met2 ;
        RECT 174.340 4434.390 200.000 4458.290 ;
      LAYER met2 ;
        RECT 4.925 4408.675 197.965 4434.110 ;
      LAYER met2 ;
        RECT 200.650 4422.195 200.930 4422.565 ;
      LAYER met2 ;
        RECT 4.925 4384.265 197.665 4408.675 ;
      LAYER met2 ;
        RECT 197.945 4384.495 200.000 4408.395 ;
        RECT 200.720 4385.165 200.860 4422.195 ;
        RECT 200.650 4384.795 200.930 4385.165 ;
        RECT 210.770 4384.795 211.050 4385.165 ;
        RECT 210.840 4347.230 210.980 4384.795 ;
        RECT 210.780 4346.910 211.040 4347.230 ;
        RECT 211.300 3871.570 211.440 4950.410 ;
        RECT 224.180 4623.165 224.320 4952.110 ;
        RECT 224.580 4951.430 224.840 4951.750 ;
        RECT 223.190 4622.795 223.470 4623.165 ;
        RECT 224.110 4622.795 224.390 4623.165 ;
        RECT 222.280 4574.370 222.540 4574.690 ;
        RECT 222.340 4443.790 222.480 4574.370 ;
        RECT 223.260 4526.605 223.400 4622.795 ;
        RECT 224.640 4622.370 224.780 4951.430 ;
        RECT 317.560 4951.070 317.700 4952.110 ;
        RECT 386.490 4951.235 386.770 4951.605 ;
        RECT 386.500 4951.090 386.760 4951.235 ;
        RECT 412.320 4951.070 412.460 4952.110 ;
        RECT 530.940 4951.770 531.200 4952.090 ;
        RECT 414.090 4951.235 414.370 4951.605 ;
        RECT 317.500 4950.750 317.760 4951.070 ;
        RECT 412.260 4950.750 412.520 4951.070 ;
        RECT 414.160 4950.730 414.300 4951.235 ;
        RECT 414.100 4950.410 414.360 4950.730 ;
        RECT 510.690 4950.555 510.970 4950.925 ;
        RECT 531.000 4950.730 531.140 4951.770 ;
        RECT 663.020 4951.410 663.160 4952.710 ;
        RECT 662.960 4951.090 663.220 4951.410 ;
        RECT 684.640 4951.070 684.780 4953.810 ;
        RECT 737.080 4952.770 737.220 4977.035 ;
        RECT 1228.300 4960.270 1228.560 4960.590 ;
        RECT 1226.000 4953.810 1226.260 4954.130 ;
        RECT 1089.840 4953.130 1090.100 4953.450 ;
        RECT 737.020 4952.450 737.280 4952.770 ;
        RECT 772.960 4952.710 773.560 4952.850 ;
        RECT 510.700 4950.410 510.960 4950.555 ;
        RECT 530.940 4950.410 531.200 4950.730 ;
        RECT 531.390 4950.555 531.670 4950.925 ;
        RECT 684.580 4950.750 684.840 4951.070 ;
        RECT 737.080 4950.730 737.220 4952.450 ;
        RECT 772.960 4952.430 773.100 4952.710 ;
        RECT 772.900 4952.110 773.160 4952.430 ;
        RECT 758.640 4951.770 758.900 4952.090 ;
        RECT 758.700 4951.410 758.840 4951.770 ;
        RECT 758.640 4951.090 758.900 4951.410 ;
        RECT 773.420 4951.070 773.560 4952.710 ;
        RECT 966.090 4951.235 966.370 4951.605 ;
        RECT 1089.900 4951.410 1090.040 4953.130 ;
        RECT 1226.060 4952.430 1226.200 4953.810 ;
        RECT 1226.000 4952.110 1226.260 4952.430 ;
        RECT 1179.540 4951.770 1179.800 4952.090 ;
        RECT 1227.840 4951.770 1228.100 4952.090 ;
        RECT 966.100 4951.090 966.360 4951.235 ;
        RECT 1089.840 4951.090 1090.100 4951.410 ;
        RECT 1091.210 4951.235 1091.490 4951.605 ;
        RECT 773.360 4950.750 773.620 4951.070 ;
        RECT 1091.280 4950.730 1091.420 4951.235 ;
        RECT 1179.600 4950.730 1179.740 4951.770 ;
        RECT 1226.980 4951.410 1227.580 4951.490 ;
        RECT 1226.980 4951.350 1227.640 4951.410 ;
        RECT 1226.980 4951.070 1227.120 4951.350 ;
        RECT 1227.380 4951.090 1227.640 4951.350 ;
        RECT 1227.900 4951.070 1228.040 4951.770 ;
        RECT 1228.360 4951.410 1228.500 4960.270 ;
        RECT 1229.740 4952.430 1229.880 4977.035 ;
        RECT 1251.760 4976.930 1252.020 4977.190 ;
        RECT 1266.465 4977.035 1266.745 4979.435 ;
        RECT 1272.905 4977.035 1273.185 4979.435 ;
        RECT 1275.665 4977.035 1275.945 4979.435 ;
        RECT 1282.105 4977.035 1282.385 4979.435 ;
        RECT 1284.865 4977.035 1285.145 4979.435 ;
        RECT 1291.305 4977.330 1291.585 4979.435 ;
        RECT 1290.920 4977.250 1291.585 4977.330 ;
        RECT 1290.860 4977.190 1291.585 4977.250 ;
        RECT 1282.180 4960.590 1282.320 4977.035 ;
        RECT 1290.860 4976.930 1291.120 4977.190 ;
        RECT 1291.305 4977.035 1291.585 4977.190 ;
        RECT 1282.120 4960.270 1282.380 4960.590 ;
        RECT 1282.180 4952.770 1282.320 4960.270 ;
        RECT 1282.120 4952.450 1282.380 4952.770 ;
        RECT 1435.290 4952.595 1435.570 4952.965 ;
        RECT 1450.010 4952.595 1450.290 4952.965 ;
        RECT 1435.300 4952.450 1435.560 4952.595 ;
        RECT 1229.680 4952.110 1229.940 4952.430 ;
        RECT 1448.640 4952.170 1448.900 4952.430 ;
        RECT 1449.560 4952.170 1449.820 4952.430 ;
        RECT 1448.640 4952.110 1449.820 4952.170 ;
        RECT 1448.700 4952.030 1449.760 4952.110 ;
        RECT 1450.080 4952.090 1450.220 4952.595 ;
        RECT 1545.240 4952.450 1545.500 4952.770 ;
        RECT 1545.300 4952.090 1545.440 4952.450 ;
        RECT 1450.020 4951.770 1450.280 4952.090 ;
        RECT 1545.240 4951.770 1545.500 4952.090 ;
        RECT 1620.280 4951.605 1620.420 4982.515 ;
      LAYER met2 ;
        RECT 1758.210 4979.715 1837.915 5188.000 ;
        RECT 1758.210 4979.435 1759.205 4979.715 ;
        RECT 1760.045 4979.435 1761.965 4979.715 ;
        RECT 1762.805 4979.435 1765.185 4979.715 ;
        RECT 1766.025 4979.435 1768.405 4979.715 ;
        RECT 1769.245 4979.435 1771.165 4979.715 ;
        RECT 1772.005 4979.435 1774.385 4979.715 ;
        RECT 1775.225 4979.435 1777.605 4979.715 ;
        RECT 1778.445 4979.435 1780.365 4979.715 ;
        RECT 1781.205 4979.435 1783.585 4979.715 ;
        RECT 1784.425 4979.435 1786.805 4979.715 ;
        RECT 1787.645 4979.435 1789.565 4979.715 ;
        RECT 1790.405 4979.435 1792.785 4979.715 ;
        RECT 1793.625 4979.435 1796.005 4979.715 ;
        RECT 1796.845 4979.435 1799.225 4979.715 ;
        RECT 1800.065 4979.435 1801.985 4979.715 ;
        RECT 1802.825 4979.435 1805.205 4979.715 ;
        RECT 1806.045 4979.435 1808.425 4979.715 ;
        RECT 1809.265 4979.435 1811.185 4979.715 ;
        RECT 1812.025 4979.435 1814.405 4979.715 ;
        RECT 1815.245 4979.435 1817.625 4979.715 ;
        RECT 1818.465 4979.435 1820.385 4979.715 ;
        RECT 1821.225 4979.435 1823.605 4979.715 ;
        RECT 1824.445 4979.435 1826.825 4979.715 ;
        RECT 1827.665 4979.435 1829.585 4979.715 ;
        RECT 1830.425 4979.435 1832.805 4979.715 ;
        RECT 1833.645 4979.435 1836.025 4979.715 ;
        RECT 1836.865 4979.435 1837.915 4979.715 ;
        RECT 2303.210 4979.715 2382.915 5188.000 ;
        RECT 2848.265 5013.940 2922.290 5183.075 ;
        RECT 2848.265 4990.335 2898.110 5013.940 ;
      LAYER met2 ;
        RECT 2848.495 4988.000 2872.395 4990.055 ;
      LAYER met2 ;
        RECT 2872.675 4990.035 2898.110 4990.335 ;
      LAYER met2 ;
        RECT 2898.390 4988.000 2922.290 5013.660 ;
        RECT 2870.030 4985.235 2870.310 4985.605 ;
      LAYER met2 ;
        RECT 2303.210 4979.435 2304.205 4979.715 ;
        RECT 2305.045 4979.435 2306.965 4979.715 ;
        RECT 2307.805 4979.435 2310.185 4979.715 ;
        RECT 2311.025 4979.435 2313.405 4979.715 ;
        RECT 2314.245 4979.435 2316.165 4979.715 ;
        RECT 2317.005 4979.435 2319.385 4979.715 ;
        RECT 2320.225 4979.435 2322.605 4979.715 ;
        RECT 2323.445 4979.435 2325.365 4979.715 ;
        RECT 2326.205 4979.435 2328.585 4979.715 ;
        RECT 2329.425 4979.435 2331.805 4979.715 ;
        RECT 2332.645 4979.435 2334.565 4979.715 ;
        RECT 2335.405 4979.435 2337.785 4979.715 ;
        RECT 2338.625 4979.435 2341.005 4979.715 ;
        RECT 2341.845 4979.435 2344.225 4979.715 ;
        RECT 2345.065 4979.435 2346.985 4979.715 ;
        RECT 2347.825 4979.435 2350.205 4979.715 ;
        RECT 2351.045 4979.435 2353.425 4979.715 ;
        RECT 2354.265 4979.435 2356.185 4979.715 ;
        RECT 2357.025 4979.435 2359.405 4979.715 ;
        RECT 2360.245 4979.435 2362.625 4979.715 ;
        RECT 2363.465 4979.435 2365.385 4979.715 ;
        RECT 2366.225 4979.435 2368.605 4979.715 ;
        RECT 2369.445 4979.435 2371.825 4979.715 ;
        RECT 2372.665 4979.435 2374.585 4979.715 ;
        RECT 2375.425 4979.435 2377.805 4979.715 ;
        RECT 2378.645 4979.435 2381.025 4979.715 ;
        RECT 2381.865 4979.435 2382.915 4979.715 ;
      LAYER met2 ;
        RECT 1759.485 4977.035 1759.765 4979.435 ;
        RECT 1774.665 4977.260 1774.945 4979.435 ;
        RECT 1796.285 4977.260 1796.565 4979.435 ;
        RECT 1774.665 4977.035 1774.980 4977.260 ;
        RECT 1796.285 4977.035 1796.600 4977.260 ;
        RECT 1811.465 4977.035 1811.745 4979.435 ;
        RECT 1817.905 4977.035 1818.185 4979.435 ;
        RECT 1820.665 4977.035 1820.945 4979.435 ;
        RECT 1827.105 4977.260 1827.385 4979.435 ;
        RECT 1827.105 4977.035 1827.420 4977.260 ;
        RECT 1829.865 4977.035 1830.145 4979.435 ;
        RECT 1836.305 4977.260 1836.585 4979.435 ;
        RECT 1836.305 4977.035 1836.620 4977.260 ;
        RECT 2304.485 4977.035 2304.765 4979.435 ;
        RECT 2319.665 4977.330 2319.945 4979.435 ;
        RECT 2341.285 4977.330 2341.565 4979.435 ;
        RECT 2341.960 4977.330 2342.220 4977.590 ;
        RECT 2319.665 4977.035 2320.080 4977.330 ;
        RECT 2341.285 4977.270 2342.220 4977.330 ;
        RECT 2341.285 4977.190 2342.160 4977.270 ;
        RECT 2341.285 4977.035 2341.565 4977.190 ;
        RECT 2356.465 4977.035 2356.745 4979.435 ;
        RECT 2362.905 4977.035 2363.185 4979.435 ;
        RECT 2365.665 4977.035 2365.945 4979.435 ;
        RECT 2372.105 4977.330 2372.385 4979.435 ;
        RECT 2372.105 4977.035 2372.520 4977.330 ;
        RECT 2374.865 4977.035 2375.145 4979.435 ;
        RECT 2380.600 4977.330 2380.860 4977.590 ;
        RECT 2381.305 4977.330 2381.585 4979.435 ;
        RECT 2380.600 4977.270 2381.585 4977.330 ;
        RECT 2380.660 4977.190 2381.585 4977.270 ;
        RECT 2381.305 4977.035 2381.585 4977.190 ;
        RECT 1628.500 4952.450 1628.760 4952.770 ;
        RECT 1628.950 4952.595 1629.230 4952.965 ;
        RECT 1738.430 4952.595 1738.710 4952.965 ;
        RECT 1628.560 4952.170 1628.700 4952.450 ;
        RECT 1629.020 4952.170 1629.160 4952.595 ;
        RECT 1738.440 4952.450 1738.700 4952.595 ;
        RECT 1774.840 4952.430 1774.980 4977.035 ;
        RECT 1796.460 4954.130 1796.600 4977.035 ;
        RECT 1796.400 4953.810 1796.660 4954.130 ;
        RECT 1827.280 4953.790 1827.420 4977.035 ;
        RECT 1836.480 4954.130 1836.620 4977.035 ;
        RECT 1836.420 4953.810 1836.680 4954.130 ;
        RECT 2319.940 4953.790 2320.080 4977.035 ;
        RECT 2372.380 4954.130 2372.520 4977.035 ;
        RECT 2370.020 4953.810 2370.280 4954.130 ;
        RECT 2372.320 4953.810 2372.580 4954.130 ;
        RECT 1827.220 4953.470 1827.480 4953.790 ;
        RECT 2319.880 4953.470 2320.140 4953.790 ;
        RECT 1827.280 4952.770 1827.420 4953.470 ;
        RECT 1827.220 4952.450 1827.480 4952.770 ;
        RECT 1628.560 4952.030 1629.160 4952.170 ;
        RECT 1774.780 4952.110 1775.040 4952.430 ;
        RECT 1228.300 4951.090 1228.560 4951.410 ;
        RECT 1380.100 4951.090 1380.360 4951.410 ;
        RECT 1474.850 4951.235 1475.130 4951.605 ;
        RECT 1620.210 4951.235 1620.490 4951.605 ;
        RECT 1474.860 4951.090 1475.120 4951.235 ;
        RECT 1226.920 4950.750 1227.180 4951.070 ;
        RECT 1227.840 4950.750 1228.100 4951.070 ;
        RECT 1379.640 4950.810 1379.900 4951.070 ;
        RECT 1380.160 4950.810 1380.300 4951.090 ;
        RECT 1379.640 4950.750 1380.300 4950.810 ;
        RECT 531.400 4950.410 531.660 4950.555 ;
        RECT 737.020 4950.410 737.280 4950.730 ;
        RECT 1091.220 4950.410 1091.480 4950.730 ;
        RECT 1179.540 4950.410 1179.800 4950.730 ;
        RECT 1379.700 4950.670 1380.300 4950.750 ;
        RECT 2370.080 4950.730 2370.220 4953.810 ;
        RECT 2856.700 4953.470 2856.960 4953.790 ;
        RECT 2856.760 4951.070 2856.900 4953.470 ;
        RECT 2870.100 4951.070 2870.240 4985.235 ;
        RECT 2856.700 4950.750 2856.960 4951.070 ;
        RECT 2870.040 4950.750 2870.300 4951.070 ;
        RECT 3373.740 4950.750 3374.000 4951.070 ;
        RECT 2370.020 4950.410 2370.280 4950.730 ;
        RECT 3365.460 4950.410 3365.720 4950.730 ;
        RECT 224.180 4622.230 224.780 4622.370 ;
        RECT 224.180 4574.690 224.320 4622.230 ;
        RECT 224.120 4574.370 224.380 4574.690 ;
        RECT 223.190 4526.235 223.470 4526.605 ;
        RECT 224.110 4526.235 224.390 4526.605 ;
        RECT 222.280 4443.470 222.540 4443.790 ;
        RECT 223.660 4443.470 223.920 4443.790 ;
        RECT 223.720 4422.565 223.860 4443.470 ;
        RECT 223.650 4422.195 223.930 4422.565 ;
        RECT 224.180 4410.325 224.320 4526.235 ;
        RECT 220.890 4409.955 221.170 4410.325 ;
        RECT 224.110 4409.955 224.390 4410.325 ;
        RECT 211.240 3871.250 211.500 3871.570 ;
        RECT 212.620 3871.250 212.880 3871.570 ;
      LAYER met2 ;
        RECT 0.000 3853.865 208.565 3854.915 ;
        RECT 0.000 3853.025 208.285 3853.865 ;
      LAYER met2 ;
        RECT 208.565 3853.305 210.965 3853.585 ;
      LAYER met2 ;
        RECT 0.000 3850.645 208.565 3853.025 ;
      LAYER met2 ;
        RECT 209.000 3851.250 209.140 3853.305 ;
        RECT 209.000 3851.110 211.440 3851.250 ;
      LAYER met2 ;
        RECT 0.000 3849.805 208.285 3850.645 ;
        RECT 0.000 3847.425 208.565 3849.805 ;
        RECT 0.000 3846.585 208.285 3847.425 ;
      LAYER met2 ;
        RECT 208.565 3846.865 210.965 3847.145 ;
      LAYER met2 ;
        RECT 0.000 3844.665 208.565 3846.585 ;
      LAYER met2 ;
        RECT 208.940 3846.090 209.200 3846.410 ;
      LAYER met2 ;
        RECT 0.000 3843.825 208.285 3844.665 ;
      LAYER met2 ;
        RECT 209.000 3844.450 209.140 3846.090 ;
        RECT 208.610 3844.385 209.140 3844.450 ;
        RECT 208.565 3844.105 210.965 3844.385 ;
      LAYER met2 ;
        RECT 0.000 3841.445 208.565 3843.825 ;
        RECT 0.000 3840.605 208.285 3841.445 ;
        RECT 0.000 3838.225 208.565 3840.605 ;
        RECT 0.000 3837.385 208.285 3838.225 ;
      LAYER met2 ;
        RECT 208.565 3837.665 210.965 3837.945 ;
      LAYER met2 ;
        RECT 0.000 3835.465 208.565 3837.385 ;
        RECT 0.000 3834.625 208.285 3835.465 ;
      LAYER met2 ;
        RECT 208.565 3834.905 210.965 3835.185 ;
      LAYER met2 ;
        RECT 0.000 3832.245 208.565 3834.625 ;
        RECT 0.000 3831.405 208.285 3832.245 ;
        RECT 0.000 3829.025 208.565 3831.405 ;
        RECT 0.000 3828.185 208.285 3829.025 ;
      LAYER met2 ;
        RECT 208.565 3828.465 210.965 3828.745 ;
      LAYER met2 ;
        RECT 0.000 3826.265 208.565 3828.185 ;
        RECT 0.000 3825.425 208.285 3826.265 ;
        RECT 0.000 3823.045 208.565 3825.425 ;
        RECT 0.000 3822.205 208.285 3823.045 ;
        RECT 0.000 3819.825 208.565 3822.205 ;
        RECT 0.000 3818.985 208.285 3819.825 ;
        RECT 0.000 3817.065 208.565 3818.985 ;
        RECT 0.000 3816.225 208.285 3817.065 ;
        RECT 0.000 3813.845 208.565 3816.225 ;
      LAYER met2 ;
        RECT 211.300 3813.850 211.440 3851.110 ;
        RECT 212.680 3846.410 212.820 3871.250 ;
        RECT 212.620 3846.090 212.880 3846.410 ;
        RECT 212.680 3836.890 212.820 3846.090 ;
        RECT 211.700 3836.570 211.960 3836.890 ;
        RECT 212.620 3836.570 212.880 3836.890 ;
      LAYER met2 ;
        RECT 0.000 3813.005 208.285 3813.845 ;
      LAYER met2 ;
        RECT 209.000 3813.710 211.440 3813.850 ;
        RECT 209.000 3813.565 209.140 3813.710 ;
        RECT 208.565 3813.285 210.965 3813.565 ;
      LAYER met2 ;
        RECT 0.000 3810.625 208.565 3813.005 ;
        RECT 0.000 3809.785 208.285 3810.625 ;
        RECT 0.000 3807.405 208.565 3809.785 ;
        RECT 0.000 3806.565 208.285 3807.405 ;
        RECT 0.000 3804.645 208.565 3806.565 ;
        RECT 0.000 3803.805 208.285 3804.645 ;
        RECT 0.000 3801.425 208.565 3803.805 ;
        RECT 0.000 3800.585 208.285 3801.425 ;
        RECT 0.000 3798.205 208.565 3800.585 ;
        RECT 0.000 3797.365 208.285 3798.205 ;
        RECT 0.000 3795.445 208.565 3797.365 ;
        RECT 0.000 3794.605 208.285 3795.445 ;
        RECT 0.000 3792.225 208.565 3794.605 ;
      LAYER met2 ;
        RECT 208.940 3792.370 209.200 3792.690 ;
      LAYER met2 ;
        RECT 0.000 3791.385 208.285 3792.225 ;
      LAYER met2 ;
        RECT 209.000 3791.945 209.140 3792.370 ;
        RECT 208.565 3791.665 210.965 3791.945 ;
      LAYER met2 ;
        RECT 0.000 3789.005 208.565 3791.385 ;
        RECT 0.000 3788.165 208.285 3789.005 ;
        RECT 0.000 3786.245 208.565 3788.165 ;
      LAYER met2 ;
        RECT 211.760 3788.010 211.900 3836.570 ;
        RECT 220.960 3792.690 221.100 4409.955 ;
        RECT 3365.520 4400.270 3365.660 4950.410 ;
        RECT 3373.800 4471.670 3373.940 4950.750 ;
        RECT 3368.680 4471.350 3368.940 4471.670 ;
        RECT 3373.740 4471.350 3374.000 4471.670 ;
        RECT 3390.300 4471.350 3390.560 4471.670 ;
        RECT 3365.460 4399.950 3365.720 4400.270 ;
        RECT 3368.220 4399.950 3368.480 4400.270 ;
        RECT 3368.280 4380.890 3368.420 4399.950 ;
        RECT 3368.220 4380.570 3368.480 4380.890 ;
        RECT 223.660 4346.910 223.920 4347.230 ;
        RECT 223.720 4278.290 223.860 4346.910 ;
        RECT 223.720 4278.150 224.320 4278.290 ;
        RECT 224.180 4250.410 224.320 4278.150 ;
        RECT 223.720 4250.270 224.320 4250.410 ;
        RECT 223.720 4181.650 223.860 4250.270 ;
        RECT 223.660 4181.330 223.920 4181.650 ;
        RECT 223.200 4180.990 223.460 4181.310 ;
        RECT 223.260 4154.110 223.400 4180.990 ;
        RECT 223.200 4153.790 223.460 4154.110 ;
        RECT 223.660 4153.790 223.920 4154.110 ;
        RECT 223.720 4058.085 223.860 4153.790 ;
        RECT 223.650 4057.715 223.930 4058.085 ;
        RECT 223.190 4057.290 223.470 4057.405 ;
        RECT 222.800 4057.150 223.470 4057.290 ;
        RECT 222.800 3988.610 222.940 4057.150 ;
        RECT 223.190 4057.035 223.470 4057.150 ;
        RECT 222.800 3988.470 223.400 3988.610 ;
        RECT 223.260 3987.930 223.400 3988.470 ;
        RECT 222.340 3987.790 223.400 3987.930 ;
        RECT 222.340 3891.970 222.480 3987.790 ;
        RECT 222.280 3891.650 222.540 3891.970 ;
        RECT 222.740 3890.970 223.000 3891.290 ;
        RECT 222.800 3794.810 222.940 3890.970 ;
        RECT 222.800 3794.670 223.860 3794.810 ;
        RECT 213.080 3792.370 213.340 3792.690 ;
        RECT 220.900 3792.370 221.160 3792.690 ;
        RECT 211.300 3787.870 211.900 3788.010 ;
      LAYER met2 ;
        RECT 0.000 3785.405 208.285 3786.245 ;
        RECT 0.000 3783.025 208.565 3785.405 ;
        RECT 0.000 3782.185 208.285 3783.025 ;
        RECT 0.000 3779.805 208.565 3782.185 ;
        RECT 0.000 3778.965 208.285 3779.805 ;
        RECT 0.000 3777.045 208.565 3778.965 ;
        RECT 0.000 3776.205 208.285 3777.045 ;
      LAYER met2 ;
        RECT 208.565 3776.485 210.965 3776.765 ;
      LAYER met2 ;
        RECT 0.000 3775.210 208.565 3776.205 ;
      LAYER met2 ;
        RECT 211.300 3254.810 211.440 3787.870 ;
        RECT 213.140 3758.010 213.280 3792.370 ;
        RECT 211.700 3757.690 211.960 3758.010 ;
        RECT 213.080 3757.690 213.340 3758.010 ;
        RECT 211.240 3254.490 211.500 3254.810 ;
      LAYER met2 ;
        RECT 0.000 3245.865 208.565 3246.915 ;
        RECT 0.000 3245.025 208.285 3245.865 ;
      LAYER met2 ;
        RECT 208.565 3245.445 210.965 3245.585 ;
        RECT 208.540 3245.370 210.965 3245.445 ;
        RECT 208.540 3245.230 211.440 3245.370 ;
      LAYER met2 ;
        RECT 0.000 3242.645 208.565 3245.025 ;
        RECT 0.000 3241.805 208.285 3242.645 ;
        RECT 0.000 3239.425 208.565 3241.805 ;
        RECT 0.000 3238.585 208.285 3239.425 ;
      LAYER met2 ;
        RECT 208.565 3238.865 210.965 3239.145 ;
      LAYER met2 ;
        RECT 0.000 3236.665 208.565 3238.585 ;
      LAYER met2 ;
        RECT 208.940 3238.170 209.200 3238.490 ;
      LAYER met2 ;
        RECT 0.000 3235.825 208.285 3236.665 ;
      LAYER met2 ;
        RECT 209.000 3236.385 209.140 3238.170 ;
        RECT 208.565 3236.105 210.965 3236.385 ;
      LAYER met2 ;
        RECT 0.000 3233.445 208.565 3235.825 ;
        RECT 0.000 3232.605 208.285 3233.445 ;
        RECT 0.000 3230.225 208.565 3232.605 ;
        RECT 0.000 3229.385 208.285 3230.225 ;
      LAYER met2 ;
        RECT 208.565 3229.665 210.965 3229.945 ;
      LAYER met2 ;
        RECT 0.000 3227.465 208.565 3229.385 ;
        RECT 0.000 3226.625 208.285 3227.465 ;
      LAYER met2 ;
        RECT 208.565 3226.905 210.965 3227.185 ;
      LAYER met2 ;
        RECT 0.000 3224.245 208.565 3226.625 ;
        RECT 0.000 3223.405 208.285 3224.245 ;
        RECT 0.000 3221.025 208.565 3223.405 ;
        RECT 0.000 3220.185 208.285 3221.025 ;
      LAYER met2 ;
        RECT 208.565 3220.465 210.965 3220.745 ;
      LAYER met2 ;
        RECT 0.000 3218.265 208.565 3220.185 ;
        RECT 0.000 3217.425 208.285 3218.265 ;
        RECT 0.000 3215.045 208.565 3217.425 ;
        RECT 0.000 3214.205 208.285 3215.045 ;
        RECT 0.000 3211.825 208.565 3214.205 ;
        RECT 0.000 3210.985 208.285 3211.825 ;
        RECT 0.000 3209.065 208.565 3210.985 ;
        RECT 0.000 3208.225 208.285 3209.065 ;
        RECT 0.000 3205.845 208.565 3208.225 ;
      LAYER met2 ;
        RECT 211.300 3205.930 211.440 3245.230 ;
      LAYER met2 ;
        RECT 0.000 3205.005 208.285 3205.845 ;
      LAYER met2 ;
        RECT 209.460 3205.790 211.440 3205.930 ;
        RECT 209.460 3205.565 209.600 3205.790 ;
        RECT 208.565 3205.285 210.965 3205.565 ;
      LAYER met2 ;
        RECT 0.000 3202.625 208.565 3205.005 ;
        RECT 0.000 3201.785 208.285 3202.625 ;
        RECT 0.000 3199.405 208.565 3201.785 ;
        RECT 0.000 3198.565 208.285 3199.405 ;
        RECT 0.000 3196.645 208.565 3198.565 ;
        RECT 0.000 3195.805 208.285 3196.645 ;
        RECT 0.000 3193.425 208.565 3195.805 ;
        RECT 0.000 3192.585 208.285 3193.425 ;
        RECT 0.000 3190.205 208.565 3192.585 ;
        RECT 0.000 3189.365 208.285 3190.205 ;
        RECT 0.000 3187.445 208.565 3189.365 ;
        RECT 0.000 3186.605 208.285 3187.445 ;
        RECT 0.000 3184.225 208.565 3186.605 ;
      LAYER met2 ;
        RECT 211.760 3186.210 211.900 3757.690 ;
        RECT 223.720 3698.850 223.860 3794.670 ;
        RECT 3368.280 3779.770 3368.420 4380.570 ;
        RECT 3368.740 3836.890 3368.880 4471.350 ;
        RECT 3390.360 4454.500 3390.500 4471.350 ;
        RECT 3390.000 4434.505 3391.485 4454.500 ;
      LAYER met2 ;
        RECT 3391.765 4434.225 3584.430 4454.510 ;
        RECT 3390.035 4420.840 3584.430 4434.225 ;
      LAYER met2 ;
        RECT 3390.000 4410.890 3390.325 4420.560 ;
        RECT 3388.520 4410.750 3390.325 4410.890 ;
        RECT 3388.520 4374.770 3388.660 4410.750 ;
        RECT 3390.000 4410.560 3390.325 4410.750 ;
      LAYER met2 ;
        RECT 3390.605 4410.280 3584.430 4420.840 ;
      LAYER met2 ;
        RECT 3389.370 4405.875 3389.650 4406.245 ;
        RECT 3389.440 4381.085 3389.580 4405.875 ;
      LAYER met2 ;
        RECT 3390.035 4400.565 3584.430 4410.280 ;
      LAYER met2 ;
        RECT 3389.370 4380.715 3389.650 4381.085 ;
        RECT 3389.380 4380.570 3389.640 4380.715 ;
        RECT 3390.000 4380.300 3393.660 4400.285 ;
      LAYER met2 ;
        RECT 3393.940 4380.300 3584.430 4400.565 ;
      LAYER met2 ;
        RECT 3373.740 4374.450 3374.000 4374.770 ;
        RECT 3388.460 4374.450 3388.720 4374.770 ;
        RECT 3368.680 3836.570 3368.940 3836.890 ;
        RECT 3367.300 3779.450 3367.560 3779.770 ;
        RECT 3368.220 3779.450 3368.480 3779.770 ;
        RECT 223.660 3698.530 223.920 3698.850 ;
        RECT 224.120 3697.850 224.380 3698.170 ;
        RECT 224.180 3670.630 224.320 3697.850 ;
        RECT 223.200 3670.310 223.460 3670.630 ;
        RECT 224.120 3670.310 224.380 3670.630 ;
        RECT 223.260 3601.950 223.400 3670.310 ;
        RECT 223.200 3601.630 223.460 3601.950 ;
        RECT 224.120 3601.630 224.380 3601.950 ;
        RECT 224.180 3574.490 224.320 3601.630 ;
        RECT 224.180 3574.350 224.780 3574.490 ;
        RECT 224.640 3525.530 224.780 3574.350 ;
        RECT 224.180 3525.390 224.780 3525.530 ;
        RECT 224.180 3505.390 224.320 3525.390 ;
        RECT 224.120 3505.070 224.380 3505.390 ;
        RECT 224.120 3504.390 224.380 3504.710 ;
        RECT 224.180 3463.910 224.320 3504.390 ;
        RECT 222.280 3463.590 222.540 3463.910 ;
        RECT 224.120 3463.590 224.380 3463.910 ;
        RECT 222.340 3367.690 222.480 3463.590 ;
        RECT 222.280 3367.370 222.540 3367.690 ;
        RECT 223.660 3367.370 223.920 3367.690 ;
        RECT 223.720 3312.610 223.860 3367.370 ;
        RECT 223.660 3312.290 223.920 3312.610 ;
        RECT 223.200 3311.610 223.460 3311.930 ;
        RECT 223.260 3270.645 223.400 3311.610 ;
        RECT 223.190 3270.275 223.470 3270.645 ;
        RECT 224.110 3270.275 224.390 3270.645 ;
        RECT 212.160 3254.490 212.420 3254.810 ;
        RECT 212.220 3238.490 212.360 3254.490 ;
        RECT 212.160 3238.170 212.420 3238.490 ;
        RECT 213.080 3238.170 213.340 3238.490 ;
        RECT 209.000 3186.070 211.900 3186.210 ;
      LAYER met2 ;
        RECT 0.000 3183.385 208.285 3184.225 ;
      LAYER met2 ;
        RECT 209.000 3183.945 209.140 3186.070 ;
        RECT 208.565 3183.665 210.965 3183.945 ;
      LAYER met2 ;
        RECT 0.000 3181.005 208.565 3183.385 ;
        RECT 0.000 3180.165 208.285 3181.005 ;
        RECT 0.000 3178.245 208.565 3180.165 ;
        RECT 0.000 3177.405 208.285 3178.245 ;
        RECT 0.000 3175.025 208.565 3177.405 ;
        RECT 0.000 3174.185 208.285 3175.025 ;
        RECT 0.000 3171.805 208.565 3174.185 ;
        RECT 0.000 3170.965 208.285 3171.805 ;
        RECT 0.000 3169.045 208.565 3170.965 ;
        RECT 0.000 3168.205 208.285 3169.045 ;
      LAYER met2 ;
        RECT 208.565 3168.485 210.965 3168.765 ;
      LAYER met2 ;
        RECT 0.000 3167.210 208.565 3168.205 ;
      LAYER met2 ;
        RECT 213.140 3118.470 213.280 3238.170 ;
        RECT 211.240 3118.150 211.500 3118.470 ;
        RECT 213.080 3118.150 213.340 3118.470 ;
        RECT 211.300 2683.690 211.440 3118.150 ;
        RECT 224.180 3092.290 224.320 3270.275 ;
        RECT 3367.360 3171.850 3367.500 3779.450 ;
        RECT 3368.740 3228.970 3368.880 3836.570 ;
        RECT 3368.680 3228.650 3368.940 3228.970 ;
        RECT 3367.300 3171.530 3367.560 3171.850 ;
        RECT 224.120 3091.970 224.380 3092.290 ;
        RECT 224.120 3091.290 224.380 3091.610 ;
        RECT 224.180 3022.590 224.320 3091.290 ;
        RECT 224.120 3022.270 224.380 3022.590 ;
        RECT 223.660 3021.930 223.920 3022.250 ;
        RECT 223.720 2925.770 223.860 3021.930 ;
        RECT 222.800 2925.630 223.860 2925.770 ;
        RECT 222.800 2898.150 222.940 2925.630 ;
        RECT 221.820 2897.830 222.080 2898.150 ;
        RECT 222.740 2897.830 223.000 2898.150 ;
        RECT 221.880 2801.590 222.020 2897.830 ;
        RECT 221.820 2801.270 222.080 2801.590 ;
        RECT 223.200 2801.270 223.460 2801.590 ;
        RECT 223.260 2732.650 223.400 2801.270 ;
        RECT 223.260 2732.510 224.320 2732.650 ;
        RECT 211.300 2683.550 213.280 2683.690 ;
      LAYER met2 ;
        RECT 0.000 2636.865 208.565 2637.915 ;
        RECT 0.000 2636.025 208.285 2636.865 ;
      LAYER met2 ;
        RECT 208.470 2636.585 208.750 2636.630 ;
        RECT 208.470 2636.305 210.965 2636.585 ;
        RECT 208.470 2636.260 208.750 2636.305 ;
        RECT 211.230 2636.260 211.510 2636.630 ;
      LAYER met2 ;
        RECT 0.000 2633.645 208.565 2636.025 ;
        RECT 0.000 2632.805 208.285 2633.645 ;
        RECT 0.000 2630.425 208.565 2632.805 ;
      LAYER met2 ;
        RECT 211.300 2632.010 211.440 2636.260 ;
        RECT 210.840 2631.870 211.440 2632.010 ;
        RECT 210.840 2630.650 210.980 2631.870 ;
        RECT 210.840 2630.510 211.900 2630.650 ;
      LAYER met2 ;
        RECT 0.000 2629.585 208.285 2630.425 ;
      LAYER met2 ;
        RECT 208.565 2629.865 210.965 2630.145 ;
      LAYER met2 ;
        RECT 0.000 2627.665 208.565 2629.585 ;
      LAYER met2 ;
        RECT 208.940 2629.230 209.200 2629.550 ;
      LAYER met2 ;
        RECT 0.000 2626.825 208.285 2627.665 ;
      LAYER met2 ;
        RECT 209.000 2627.385 209.140 2629.230 ;
        RECT 208.565 2627.105 210.965 2627.385 ;
      LAYER met2 ;
        RECT 0.000 2624.445 208.565 2626.825 ;
        RECT 0.000 2623.605 208.285 2624.445 ;
        RECT 0.000 2621.225 208.565 2623.605 ;
        RECT 0.000 2620.385 208.285 2621.225 ;
      LAYER met2 ;
        RECT 208.565 2620.665 210.965 2620.945 ;
      LAYER met2 ;
        RECT 0.000 2618.465 208.565 2620.385 ;
        RECT 0.000 2617.625 208.285 2618.465 ;
      LAYER met2 ;
        RECT 208.565 2617.905 210.965 2618.185 ;
      LAYER met2 ;
        RECT 0.000 2615.245 208.565 2617.625 ;
        RECT 0.000 2614.405 208.285 2615.245 ;
        RECT 0.000 2612.025 208.565 2614.405 ;
        RECT 0.000 2611.185 208.285 2612.025 ;
      LAYER met2 ;
        RECT 208.565 2611.465 210.965 2611.745 ;
      LAYER met2 ;
        RECT 0.000 2609.265 208.565 2611.185 ;
        RECT 0.000 2608.425 208.285 2609.265 ;
        RECT 0.000 2606.045 208.565 2608.425 ;
        RECT 0.000 2605.205 208.285 2606.045 ;
        RECT 0.000 2602.825 208.565 2605.205 ;
        RECT 0.000 2601.985 208.285 2602.825 ;
        RECT 0.000 2600.065 208.565 2601.985 ;
        RECT 0.000 2599.225 208.285 2600.065 ;
        RECT 0.000 2596.845 208.565 2599.225 ;
        RECT 0.000 2596.005 208.285 2596.845 ;
      LAYER met2 ;
        RECT 211.760 2596.650 211.900 2630.510 ;
        RECT 213.140 2629.550 213.280 2683.550 ;
        RECT 213.080 2629.230 213.340 2629.550 ;
        RECT 224.180 2608.470 224.320 2732.510 ;
        RECT 3368.740 2614.590 3368.880 3228.650 ;
        RECT 3369.140 3171.530 3369.400 3171.850 ;
        RECT 3369.200 2636.350 3369.340 3171.530 ;
        RECT 3369.140 2636.030 3369.400 2636.350 ;
        RECT 3369.140 2635.350 3369.400 2635.670 ;
        RECT 3367.300 2614.270 3367.560 2614.590 ;
        RECT 3368.680 2614.270 3368.940 2614.590 ;
        RECT 223.660 2608.150 223.920 2608.470 ;
        RECT 224.120 2608.150 224.380 2608.470 ;
        RECT 209.460 2596.565 211.900 2596.650 ;
        RECT 208.565 2596.510 211.900 2596.565 ;
        RECT 208.565 2596.285 210.965 2596.510 ;
      LAYER met2 ;
        RECT 0.000 2593.625 208.565 2596.005 ;
        RECT 0.000 2592.785 208.285 2593.625 ;
        RECT 0.000 2590.405 208.565 2592.785 ;
        RECT 0.000 2589.565 208.285 2590.405 ;
        RECT 0.000 2587.645 208.565 2589.565 ;
        RECT 0.000 2586.805 208.285 2587.645 ;
        RECT 0.000 2584.425 208.565 2586.805 ;
        RECT 0.000 2583.585 208.285 2584.425 ;
        RECT 0.000 2581.205 208.565 2583.585 ;
        RECT 0.000 2580.365 208.285 2581.205 ;
        RECT 0.000 2578.445 208.565 2580.365 ;
        RECT 0.000 2577.605 208.285 2578.445 ;
        RECT 0.000 2575.225 208.565 2577.605 ;
        RECT 0.000 2574.385 208.285 2575.225 ;
      LAYER met2 ;
        RECT 208.565 2574.890 210.965 2574.945 ;
        RECT 208.565 2574.750 212.360 2574.890 ;
        RECT 208.565 2574.665 210.965 2574.750 ;
      LAYER met2 ;
        RECT 0.000 2572.005 208.565 2574.385 ;
        RECT 0.000 2571.165 208.285 2572.005 ;
        RECT 0.000 2569.245 208.565 2571.165 ;
        RECT 0.000 2568.405 208.285 2569.245 ;
        RECT 0.000 2566.025 208.565 2568.405 ;
        RECT 0.000 2565.185 208.285 2566.025 ;
        RECT 0.000 2562.805 208.565 2565.185 ;
        RECT 0.000 2561.965 208.285 2562.805 ;
        RECT 0.000 2560.045 208.565 2561.965 ;
        RECT 0.000 2559.205 208.285 2560.045 ;
      LAYER met2 ;
        RECT 208.565 2559.485 210.965 2559.765 ;
      LAYER met2 ;
        RECT 0.000 2558.210 208.565 2559.205 ;
        RECT 0.000 2027.865 208.565 2028.915 ;
        RECT 0.000 2027.025 208.285 2027.865 ;
      LAYER met2 ;
        RECT 208.565 2027.490 210.965 2027.585 ;
        RECT 208.565 2027.350 211.440 2027.490 ;
        RECT 208.565 2027.305 210.965 2027.350 ;
      LAYER met2 ;
        RECT 0.000 2024.645 208.565 2027.025 ;
        RECT 0.000 2023.805 208.285 2024.645 ;
        RECT 0.000 2021.425 208.565 2023.805 ;
        RECT 0.000 2020.585 208.285 2021.425 ;
      LAYER met2 ;
        RECT 208.565 2020.865 210.965 2021.145 ;
      LAYER met2 ;
        RECT 0.000 2018.665 208.565 2020.585 ;
        RECT 0.000 2017.825 208.285 2018.665 ;
      LAYER met2 ;
        RECT 208.565 2018.105 210.965 2018.385 ;
      LAYER met2 ;
        RECT 0.000 2015.445 208.565 2017.825 ;
      LAYER met2 ;
        RECT 209.000 2015.850 209.140 2018.105 ;
        RECT 208.940 2015.530 209.200 2015.850 ;
      LAYER met2 ;
        RECT 0.000 2014.605 208.285 2015.445 ;
        RECT 0.000 2012.225 208.565 2014.605 ;
        RECT 0.000 2011.385 208.285 2012.225 ;
      LAYER met2 ;
        RECT 208.565 2011.665 210.965 2011.945 ;
      LAYER met2 ;
        RECT 0.000 2009.465 208.565 2011.385 ;
        RECT 0.000 2008.625 208.285 2009.465 ;
      LAYER met2 ;
        RECT 208.565 2008.905 210.965 2009.185 ;
      LAYER met2 ;
        RECT 0.000 2006.245 208.565 2008.625 ;
        RECT 0.000 2005.405 208.285 2006.245 ;
        RECT 0.000 2003.025 208.565 2005.405 ;
        RECT 0.000 2002.185 208.285 2003.025 ;
      LAYER met2 ;
        RECT 208.565 2002.465 210.965 2002.745 ;
      LAYER met2 ;
        RECT 0.000 2000.265 208.565 2002.185 ;
        RECT 0.000 1999.425 208.285 2000.265 ;
        RECT 0.000 1997.045 208.565 1999.425 ;
        RECT 0.000 1996.205 208.285 1997.045 ;
        RECT 0.000 1993.825 208.565 1996.205 ;
        RECT 0.000 1992.985 208.285 1993.825 ;
        RECT 0.000 1991.065 208.565 1992.985 ;
        RECT 0.000 1990.225 208.285 1991.065 ;
        RECT 0.000 1987.845 208.565 1990.225 ;
      LAYER met2 ;
        RECT 211.300 1988.050 211.440 2027.350 ;
        RECT 209.000 1987.910 211.440 1988.050 ;
      LAYER met2 ;
        RECT 0.000 1987.005 208.285 1987.845 ;
      LAYER met2 ;
        RECT 209.000 1987.565 209.140 1987.910 ;
        RECT 208.565 1987.285 210.965 1987.565 ;
        RECT 208.610 1987.230 209.140 1987.285 ;
      LAYER met2 ;
        RECT 0.000 1984.625 208.565 1987.005 ;
        RECT 0.000 1983.785 208.285 1984.625 ;
        RECT 0.000 1981.405 208.565 1983.785 ;
        RECT 0.000 1980.565 208.285 1981.405 ;
        RECT 0.000 1978.645 208.565 1980.565 ;
        RECT 0.000 1977.805 208.285 1978.645 ;
        RECT 0.000 1975.425 208.565 1977.805 ;
        RECT 0.000 1974.585 208.285 1975.425 ;
        RECT 0.000 1972.205 208.565 1974.585 ;
        RECT 0.000 1971.365 208.285 1972.205 ;
        RECT 0.000 1969.445 208.565 1971.365 ;
        RECT 0.000 1968.605 208.285 1969.445 ;
        RECT 0.000 1966.225 208.565 1968.605 ;
      LAYER met2 ;
        RECT 212.220 1968.590 212.360 2574.750 ;
        RECT 223.720 2521.430 223.860 2608.150 ;
        RECT 222.740 2521.110 223.000 2521.430 ;
        RECT 223.660 2521.110 223.920 2521.430 ;
        RECT 222.800 2442.550 222.940 2521.110 ;
        RECT 222.740 2442.230 223.000 2442.550 ;
        RECT 223.660 2442.230 223.920 2442.550 ;
        RECT 223.720 2346.670 223.860 2442.230 ;
        RECT 223.660 2346.350 223.920 2346.670 ;
        RECT 223.200 2345.670 223.460 2345.990 ;
        RECT 223.260 2318.450 223.400 2345.670 ;
        RECT 223.200 2318.130 223.460 2318.450 ;
        RECT 224.120 2318.130 224.380 2318.450 ;
        RECT 224.180 2222.085 224.320 2318.130 ;
        RECT 223.190 2221.715 223.470 2222.085 ;
        RECT 224.110 2221.715 224.390 2222.085 ;
        RECT 223.200 2221.570 223.460 2221.715 ;
        RECT 224.120 2221.570 224.380 2221.715 ;
        RECT 224.180 2152.610 224.320 2221.570 ;
        RECT 223.720 2152.470 224.320 2152.610 ;
        RECT 223.720 2056.050 223.860 2152.470 ;
        RECT 223.720 2055.910 224.780 2056.050 ;
        RECT 212.620 2015.530 212.880 2015.850 ;
        RECT 208.940 1968.270 209.200 1968.590 ;
        RECT 212.160 1968.270 212.420 1968.590 ;
      LAYER met2 ;
        RECT 0.000 1965.385 208.285 1966.225 ;
      LAYER met2 ;
        RECT 209.000 1965.945 209.140 1968.270 ;
        RECT 208.565 1965.665 210.965 1965.945 ;
      LAYER met2 ;
        RECT 0.000 1963.005 208.565 1965.385 ;
        RECT 0.000 1962.165 208.285 1963.005 ;
        RECT 0.000 1960.245 208.565 1962.165 ;
        RECT 0.000 1959.405 208.285 1960.245 ;
        RECT 0.000 1957.025 208.565 1959.405 ;
        RECT 0.000 1956.185 208.285 1957.025 ;
        RECT 0.000 1953.805 208.565 1956.185 ;
        RECT 0.000 1952.965 208.285 1953.805 ;
        RECT 0.000 1951.045 208.565 1952.965 ;
        RECT 0.000 1950.205 208.285 1951.045 ;
      LAYER met2 ;
        RECT 208.565 1950.485 210.965 1950.765 ;
      LAYER met2 ;
        RECT 0.000 1949.210 208.565 1950.205 ;
        RECT 0.000 1419.865 208.565 1420.915 ;
        RECT 0.000 1419.025 208.285 1419.865 ;
      LAYER met2 ;
        RECT 208.565 1419.570 210.965 1419.585 ;
        RECT 208.565 1419.430 211.440 1419.570 ;
        RECT 208.565 1419.305 210.965 1419.430 ;
      LAYER met2 ;
        RECT 0.000 1416.645 208.565 1419.025 ;
        RECT 0.000 1415.805 208.285 1416.645 ;
        RECT 0.000 1413.425 208.565 1415.805 ;
        RECT 0.000 1412.585 208.285 1413.425 ;
      LAYER met2 ;
        RECT 208.565 1412.865 210.965 1413.145 ;
      LAYER met2 ;
        RECT 0.000 1410.665 208.565 1412.585 ;
        RECT 0.000 1409.825 208.285 1410.665 ;
      LAYER met2 ;
        RECT 208.565 1410.105 210.965 1410.385 ;
      LAYER met2 ;
        RECT 0.000 1407.445 208.565 1409.825 ;
      LAYER met2 ;
        RECT 209.000 1407.930 209.140 1410.105 ;
        RECT 208.940 1407.610 209.200 1407.930 ;
      LAYER met2 ;
        RECT 0.000 1406.605 208.285 1407.445 ;
        RECT 0.000 1404.225 208.565 1406.605 ;
        RECT 0.000 1403.385 208.285 1404.225 ;
      LAYER met2 ;
        RECT 208.565 1403.665 210.965 1403.945 ;
      LAYER met2 ;
        RECT 0.000 1401.465 208.565 1403.385 ;
        RECT 0.000 1400.625 208.285 1401.465 ;
      LAYER met2 ;
        RECT 208.565 1400.905 210.965 1401.185 ;
      LAYER met2 ;
        RECT 0.000 1398.245 208.565 1400.625 ;
        RECT 0.000 1397.405 208.285 1398.245 ;
        RECT 0.000 1395.025 208.565 1397.405 ;
        RECT 0.000 1394.185 208.285 1395.025 ;
      LAYER met2 ;
        RECT 208.565 1394.465 210.965 1394.745 ;
      LAYER met2 ;
        RECT 0.000 1392.265 208.565 1394.185 ;
        RECT 0.000 1391.425 208.285 1392.265 ;
        RECT 0.000 1389.045 208.565 1391.425 ;
        RECT 0.000 1388.205 208.285 1389.045 ;
        RECT 0.000 1385.825 208.565 1388.205 ;
        RECT 0.000 1384.985 208.285 1385.825 ;
        RECT 0.000 1383.065 208.565 1384.985 ;
        RECT 0.000 1382.225 208.285 1383.065 ;
        RECT 0.000 1379.845 208.565 1382.225 ;
      LAYER met2 ;
        RECT 211.300 1380.130 211.440 1419.430 ;
        RECT 209.000 1379.990 211.440 1380.130 ;
      LAYER met2 ;
        RECT 0.000 1379.005 208.285 1379.845 ;
      LAYER met2 ;
        RECT 209.000 1379.565 209.140 1379.990 ;
        RECT 208.565 1379.285 210.965 1379.565 ;
      LAYER met2 ;
        RECT 0.000 1376.625 208.565 1379.005 ;
        RECT 0.000 1375.785 208.285 1376.625 ;
        RECT 0.000 1373.405 208.565 1375.785 ;
        RECT 0.000 1372.565 208.285 1373.405 ;
        RECT 0.000 1370.645 208.565 1372.565 ;
        RECT 0.000 1369.805 208.285 1370.645 ;
        RECT 0.000 1367.425 208.565 1369.805 ;
        RECT 0.000 1366.585 208.285 1367.425 ;
        RECT 0.000 1364.205 208.565 1366.585 ;
        RECT 0.000 1363.365 208.285 1364.205 ;
        RECT 0.000 1361.445 208.565 1363.365 ;
        RECT 0.000 1360.605 208.285 1361.445 ;
      LAYER met2 ;
        RECT 212.220 1360.670 212.360 1968.270 ;
        RECT 212.680 1407.930 212.820 2015.530 ;
        RECT 224.640 1979.890 224.780 2055.910 ;
        RECT 3367.360 2007.010 3367.500 2614.270 ;
        RECT 3369.200 2608.470 3369.340 2635.350 ;
        RECT 3369.140 2608.150 3369.400 2608.470 ;
        RECT 3370.060 2608.150 3370.320 2608.470 ;
        RECT 3370.120 2565.630 3370.260 2608.150 ;
        RECT 3368.220 2565.310 3368.480 2565.630 ;
        RECT 3370.060 2565.310 3370.320 2565.630 ;
        RECT 3367.300 2006.690 3367.560 2007.010 ;
        RECT 224.180 1979.750 224.780 1979.890 ;
        RECT 224.180 1960.090 224.320 1979.750 ;
        RECT 224.120 1959.770 224.380 1960.090 ;
        RECT 224.120 1959.090 224.380 1959.410 ;
        RECT 224.180 1835.650 224.320 1959.090 ;
        RECT 3368.280 1958.925 3368.420 2565.310 ;
        RECT 3369.140 2006.690 3369.400 2007.010 ;
        RECT 3368.210 1958.555 3368.490 1958.925 ;
        RECT 3368.220 1958.410 3368.480 1958.555 ;
        RECT 3368.280 1958.255 3368.420 1958.410 ;
        RECT 223.660 1835.330 223.920 1835.650 ;
        RECT 224.120 1835.330 224.380 1835.650 ;
        RECT 223.720 1835.165 223.860 1835.330 ;
        RECT 223.650 1834.795 223.930 1835.165 ;
        RECT 224.110 1765.435 224.390 1765.805 ;
        RECT 224.180 1738.750 224.320 1765.435 ;
        RECT 222.280 1738.430 222.540 1738.750 ;
        RECT 224.120 1738.430 224.380 1738.750 ;
        RECT 222.340 1642.530 222.480 1738.430 ;
        RECT 222.280 1642.210 222.540 1642.530 ;
        RECT 223.660 1642.210 223.920 1642.530 ;
        RECT 223.720 1573.510 223.860 1642.210 ;
        RECT 222.740 1573.190 223.000 1573.510 ;
        RECT 223.660 1573.190 223.920 1573.510 ;
        RECT 222.800 1545.630 222.940 1573.190 ;
        RECT 222.740 1545.310 223.000 1545.630 ;
        RECT 223.660 1545.310 223.920 1545.630 ;
        RECT 223.720 1476.610 223.860 1545.310 ;
        RECT 222.740 1476.290 223.000 1476.610 ;
        RECT 223.660 1476.290 223.920 1476.610 ;
        RECT 222.800 1449.070 222.940 1476.290 ;
        RECT 222.740 1448.750 223.000 1449.070 ;
        RECT 224.120 1448.750 224.380 1449.070 ;
        RECT 212.620 1407.610 212.880 1407.930 ;
      LAYER met2 ;
        RECT 0.000 1358.225 208.565 1360.605 ;
      LAYER met2 ;
        RECT 208.940 1360.350 209.200 1360.670 ;
        RECT 212.160 1360.350 212.420 1360.670 ;
      LAYER met2 ;
        RECT 0.000 1357.385 208.285 1358.225 ;
      LAYER met2 ;
        RECT 209.000 1357.945 209.140 1360.350 ;
        RECT 208.565 1357.665 210.965 1357.945 ;
      LAYER met2 ;
        RECT 0.000 1355.005 208.565 1357.385 ;
        RECT 0.000 1354.165 208.285 1355.005 ;
        RECT 0.000 1352.245 208.565 1354.165 ;
        RECT 0.000 1351.405 208.285 1352.245 ;
        RECT 0.000 1349.025 208.565 1351.405 ;
        RECT 0.000 1348.185 208.285 1349.025 ;
        RECT 0.000 1345.805 208.565 1348.185 ;
        RECT 0.000 1344.965 208.285 1345.805 ;
        RECT 0.000 1343.045 208.565 1344.965 ;
        RECT 0.000 1342.205 208.285 1343.045 ;
      LAYER met2 ;
        RECT 208.565 1342.485 210.965 1342.765 ;
      LAYER met2 ;
        RECT 0.000 1341.210 208.565 1342.205 ;
        RECT 0.000 810.865 208.565 811.915 ;
        RECT 0.000 810.025 208.285 810.865 ;
      LAYER met2 ;
        RECT 208.565 810.515 210.965 810.585 ;
        RECT 208.565 810.375 211.440 810.515 ;
        RECT 208.565 810.305 210.965 810.375 ;
      LAYER met2 ;
        RECT 0.000 807.645 208.565 810.025 ;
        RECT 0.000 806.805 208.285 807.645 ;
        RECT 0.000 804.425 208.565 806.805 ;
        RECT 0.000 803.585 208.285 804.425 ;
      LAYER met2 ;
        RECT 208.565 803.865 210.965 804.145 ;
      LAYER met2 ;
        RECT 0.000 801.665 208.565 803.585 ;
        RECT 0.000 800.825 208.285 801.665 ;
      LAYER met2 ;
        RECT 208.610 801.385 209.140 801.450 ;
        RECT 208.565 801.105 210.965 801.385 ;
      LAYER met2 ;
        RECT 0.000 798.445 208.565 800.825 ;
      LAYER met2 ;
        RECT 209.000 800.350 209.140 801.105 ;
        RECT 208.940 800.030 209.200 800.350 ;
      LAYER met2 ;
        RECT 0.000 797.605 208.285 798.445 ;
        RECT 0.000 795.225 208.565 797.605 ;
        RECT 0.000 794.385 208.285 795.225 ;
      LAYER met2 ;
        RECT 208.565 794.665 210.965 794.945 ;
      LAYER met2 ;
        RECT 0.000 792.465 208.565 794.385 ;
        RECT 0.000 791.625 208.285 792.465 ;
      LAYER met2 ;
        RECT 208.565 791.905 210.965 792.185 ;
      LAYER met2 ;
        RECT 0.000 789.245 208.565 791.625 ;
        RECT 0.000 788.405 208.285 789.245 ;
        RECT 0.000 786.025 208.565 788.405 ;
        RECT 0.000 785.185 208.285 786.025 ;
      LAYER met2 ;
        RECT 208.565 785.465 210.965 785.745 ;
      LAYER met2 ;
        RECT 0.000 783.265 208.565 785.185 ;
        RECT 0.000 782.425 208.285 783.265 ;
        RECT 0.000 780.045 208.565 782.425 ;
        RECT 0.000 779.205 208.285 780.045 ;
        RECT 0.000 776.825 208.565 779.205 ;
        RECT 0.000 775.985 208.285 776.825 ;
        RECT 0.000 774.065 208.565 775.985 ;
        RECT 0.000 773.225 208.285 774.065 ;
        RECT 0.000 770.845 208.565 773.225 ;
      LAYER met2 ;
        RECT 211.300 772.890 211.440 810.375 ;
        RECT 209.460 772.750 211.440 772.890 ;
      LAYER met2 ;
        RECT 0.000 770.005 208.285 770.845 ;
      LAYER met2 ;
        RECT 209.460 770.565 209.600 772.750 ;
        RECT 208.565 770.285 210.965 770.565 ;
      LAYER met2 ;
        RECT 0.000 767.625 208.565 770.005 ;
        RECT 0.000 766.785 208.285 767.625 ;
        RECT 0.000 764.405 208.565 766.785 ;
        RECT 0.000 763.565 208.285 764.405 ;
        RECT 0.000 761.645 208.565 763.565 ;
        RECT 0.000 760.805 208.285 761.645 ;
        RECT 0.000 758.425 208.565 760.805 ;
        RECT 0.000 757.585 208.285 758.425 ;
        RECT 0.000 755.205 208.565 757.585 ;
        RECT 0.000 754.365 208.285 755.205 ;
        RECT 0.000 752.445 208.565 754.365 ;
        RECT 0.000 751.605 208.285 752.445 ;
        RECT 0.000 749.225 208.565 751.605 ;
      LAYER met2 ;
        RECT 212.220 751.050 212.360 1360.350 ;
        RECT 212.680 800.350 212.820 1407.610 ;
        RECT 224.180 1379.710 224.320 1448.750 ;
        RECT 3369.200 1419.150 3369.340 2006.690 ;
        RECT 3369.590 1932.035 3369.870 1932.405 ;
        RECT 3369.660 1931.870 3369.800 1932.035 ;
        RECT 3369.600 1931.550 3369.860 1931.870 ;
        RECT 3370.060 1931.550 3370.320 1931.870 ;
        RECT 3370.120 1738.490 3370.260 1931.550 ;
        RECT 3369.660 1738.350 3370.260 1738.490 ;
        RECT 3369.660 1690.890 3369.800 1738.350 ;
        RECT 3369.660 1690.750 3370.260 1690.890 ;
        RECT 3370.120 1573.930 3370.260 1690.750 ;
        RECT 3370.120 1573.790 3370.720 1573.930 ;
        RECT 3370.580 1545.970 3370.720 1573.790 ;
        RECT 3369.600 1545.650 3369.860 1545.970 ;
        RECT 3370.520 1545.650 3370.780 1545.970 ;
        RECT 3369.660 1545.290 3369.800 1545.650 ;
        RECT 3369.600 1544.970 3369.860 1545.290 ;
        RECT 3370.520 1544.970 3370.780 1545.290 ;
        RECT 3369.140 1418.890 3369.400 1419.150 ;
        RECT 3368.280 1418.830 3369.400 1418.890 ;
        RECT 3368.280 1418.750 3369.340 1418.830 ;
        RECT 222.740 1379.390 223.000 1379.710 ;
        RECT 224.120 1379.390 224.380 1379.710 ;
        RECT 222.800 1352.510 222.940 1379.390 ;
        RECT 221.820 1352.190 222.080 1352.510 ;
        RECT 222.740 1352.190 223.000 1352.510 ;
        RECT 221.880 1256.290 222.020 1352.190 ;
        RECT 221.820 1255.970 222.080 1256.290 ;
        RECT 223.200 1255.970 223.460 1256.290 ;
        RECT 223.260 1187.010 223.400 1255.970 ;
        RECT 223.260 1186.870 224.320 1187.010 ;
        RECT 224.180 1062.830 224.320 1186.870 ;
        RECT 223.660 1062.510 223.920 1062.830 ;
        RECT 224.120 1062.510 224.380 1062.830 ;
        RECT 223.720 993.890 223.860 1062.510 ;
        RECT 223.720 993.750 224.320 993.890 ;
        RECT 224.180 966.010 224.320 993.750 ;
        RECT 223.720 965.870 224.320 966.010 ;
        RECT 223.720 897.250 223.860 965.870 ;
        RECT 223.660 896.930 223.920 897.250 ;
        RECT 223.200 896.590 223.460 896.910 ;
        RECT 223.260 869.710 223.400 896.590 ;
        RECT 223.200 869.390 223.460 869.710 ;
        RECT 223.660 869.390 223.920 869.710 ;
        RECT 212.620 800.030 212.880 800.350 ;
        RECT 208.940 750.730 209.200 751.050 ;
        RECT 212.160 750.730 212.420 751.050 ;
      LAYER met2 ;
        RECT 0.000 748.385 208.285 749.225 ;
      LAYER met2 ;
        RECT 209.000 748.945 209.140 750.730 ;
        RECT 208.565 748.665 210.965 748.945 ;
      LAYER met2 ;
        RECT 0.000 746.005 208.565 748.385 ;
        RECT 0.000 745.165 208.285 746.005 ;
        RECT 0.000 743.245 208.565 745.165 ;
        RECT 0.000 742.405 208.285 743.245 ;
        RECT 0.000 740.025 208.565 742.405 ;
        RECT 0.000 739.185 208.285 740.025 ;
        RECT 0.000 736.805 208.565 739.185 ;
        RECT 0.000 735.965 208.285 736.805 ;
        RECT 0.000 734.045 208.565 735.965 ;
        RECT 0.000 733.205 208.285 734.045 ;
      LAYER met2 ;
        RECT 208.565 733.485 210.965 733.765 ;
      LAYER met2 ;
        RECT 0.000 732.210 208.565 733.205 ;
      LAYER met2 ;
        RECT 212.220 228.470 212.360 750.730 ;
        RECT 212.160 228.150 212.420 228.470 ;
        RECT 212.680 213.850 212.820 800.030 ;
        RECT 223.720 773.685 223.860 869.390 ;
        RECT 3368.280 788.790 3368.420 1418.750 ;
        RECT 3370.580 1345.710 3370.720 1544.970 ;
        RECT 3369.140 1345.390 3369.400 1345.710 ;
        RECT 3370.520 1345.390 3370.780 1345.710 ;
        RECT 3369.200 1090.450 3369.340 1345.390 ;
        RECT 3369.200 1090.310 3369.800 1090.450 ;
        RECT 3369.660 897.250 3369.800 1090.310 ;
        RECT 3368.680 896.930 3368.940 897.250 ;
        RECT 3369.600 896.930 3369.860 897.250 ;
        RECT 3368.220 788.470 3368.480 788.790 ;
        RECT 223.650 773.315 223.930 773.685 ;
        RECT 223.190 772.890 223.470 773.005 ;
        RECT 222.800 772.750 223.470 772.890 ;
        RECT 222.800 704.210 222.940 772.750 ;
        RECT 223.190 772.635 223.470 772.750 ;
        RECT 3367.300 741.210 3367.560 741.530 ;
        RECT 222.800 704.070 223.400 704.210 ;
        RECT 223.260 703.530 223.400 704.070 ;
        RECT 222.800 703.390 223.400 703.530 ;
        RECT 222.800 615.130 222.940 703.390 ;
        RECT 222.800 614.990 223.400 615.130 ;
        RECT 223.260 580.030 223.400 614.990 ;
        RECT 223.200 579.710 223.460 580.030 ;
        RECT 223.660 578.690 223.920 579.010 ;
        RECT 223.720 434.930 223.860 578.690 ;
        RECT 223.720 434.790 224.320 434.930 ;
        RECT 224.180 387.250 224.320 434.790 ;
        RECT 224.120 386.930 224.380 387.250 ;
        RECT 224.120 386.250 224.380 386.570 ;
        RECT 224.180 386.085 224.320 386.250 ;
        RECT 224.110 385.715 224.390 386.085 ;
        RECT 224.110 290.090 224.390 290.205 ;
        RECT 224.110 289.950 224.780 290.090 ;
        RECT 224.110 289.835 224.390 289.950 ;
        RECT 224.640 227.790 224.780 289.950 ;
        RECT 2911.900 228.490 2912.160 228.810 ;
        RECT 1257.740 228.150 1258.000 228.470 ;
        RECT 2348.860 228.150 2349.120 228.470 ;
        RECT 224.580 227.470 224.840 227.790 ;
        RECT 741.160 221.690 741.420 222.010 ;
        RECT 212.620 213.530 212.880 213.850 ;
        RECT 676.290 202.115 676.570 202.485 ;
        RECT 676.360 200.000 676.500 202.115 ;
        RECT 741.220 201.125 741.360 221.690 ;
        RECT 1257.800 221.330 1257.940 228.150 ;
        RECT 1800.080 227.470 1800.340 227.790 ;
        RECT 1257.740 221.010 1258.000 221.330 ;
        RECT 1753.610 221.155 1753.890 221.525 ;
        RECT 1793.630 221.155 1793.910 221.525 ;
        RECT 741.150 200.755 741.430 201.125 ;
        RECT 1211.510 200.610 1211.770 200.930 ;
        RECT 1211.570 200.000 1211.710 200.610 ;
        RECT 1257.800 200.590 1257.940 221.010 ;
        RECT 1283.040 213.530 1283.300 213.850 ;
        RECT 1283.100 207.730 1283.240 213.530 ;
        RECT 1753.680 210.965 1753.820 221.155 ;
        RECT 1784.900 211.150 1785.160 211.470 ;
        RECT 1753.415 209.030 1753.820 210.965 ;
        RECT 1753.415 208.565 1753.695 209.030 ;
        RECT 1759.855 208.565 1760.135 210.965 ;
        RECT 1762.615 209.170 1762.895 210.965 ;
        RECT 1765.835 209.170 1766.115 210.965 ;
        RECT 1762.615 209.090 1763.480 209.170 ;
        RECT 1765.835 209.090 1766.700 209.170 ;
        RECT 1762.615 209.030 1763.540 209.090 ;
        RECT 1762.615 208.565 1762.895 209.030 ;
        RECT 1763.280 208.770 1763.540 209.030 ;
        RECT 1765.835 209.030 1766.760 209.090 ;
        RECT 1765.835 208.565 1766.115 209.030 ;
        RECT 1766.500 208.770 1766.760 209.030 ;
        RECT 1769.055 208.565 1769.335 210.965 ;
        RECT 1771.815 208.565 1772.095 210.965 ;
        RECT 1775.035 209.170 1775.315 210.965 ;
        RECT 1774.380 209.090 1775.315 209.170 ;
        RECT 1774.320 209.030 1775.315 209.090 ;
        RECT 1774.320 208.770 1774.580 209.030 ;
        RECT 1775.035 208.565 1775.315 209.030 ;
        RECT 1778.255 208.565 1778.535 210.965 ;
        RECT 1781.015 209.170 1781.295 210.965 ;
        RECT 1780.360 209.090 1781.295 209.170 ;
        RECT 1780.300 209.030 1781.295 209.090 ;
        RECT 1780.300 208.770 1780.560 209.030 ;
        RECT 1781.015 208.565 1781.295 209.030 ;
        RECT 1784.235 209.170 1784.515 210.965 ;
        RECT 1784.960 209.430 1785.100 211.150 ;
        RECT 1793.700 210.965 1793.840 221.155 ;
        RECT 1800.140 210.965 1800.280 227.470 ;
        RECT 1815.260 221.690 1815.520 222.010 ;
        RECT 1821.240 221.690 1821.500 222.010 ;
        RECT 1824.460 221.690 1824.720 222.010 ;
        RECT 2304.700 221.690 2304.960 222.010 ;
        RECT 1815.320 210.965 1815.460 221.690 ;
        RECT 1821.300 220.990 1821.440 221.690 ;
        RECT 1821.240 220.670 1821.500 220.990 ;
        RECT 1824.520 210.965 1824.660 221.690 ;
        RECT 1827.680 221.350 1827.940 221.670 ;
        RECT 1827.740 211.470 1827.880 221.350 ;
        RECT 1827.680 211.150 1827.940 211.470 ;
        RECT 1827.740 210.965 1827.880 211.150 ;
        RECT 1784.900 209.170 1785.160 209.430 ;
        RECT 1787.455 209.170 1787.735 210.965 ;
        RECT 1784.235 209.110 1785.160 209.170 ;
        RECT 1784.235 209.030 1785.100 209.110 ;
        RECT 1786.800 209.090 1787.735 209.170 ;
        RECT 1786.740 209.030 1787.735 209.090 ;
        RECT 1784.235 208.565 1784.515 209.030 ;
        RECT 1786.740 208.770 1787.000 209.030 ;
        RECT 1787.455 208.565 1787.735 209.030 ;
        RECT 1790.215 208.565 1790.495 210.965 ;
        RECT 1793.435 209.030 1793.840 210.965 ;
        RECT 1799.875 209.030 1800.280 210.965 ;
        RECT 1802.635 209.170 1802.915 210.965 ;
        RECT 1805.855 209.170 1806.135 210.965 ;
        RECT 1807.500 209.695 1808.100 209.835 ;
        RECT 1807.500 209.170 1807.640 209.695 ;
        RECT 1801.980 209.090 1807.640 209.170 ;
        RECT 1801.920 209.030 1807.640 209.090 ;
        RECT 1807.960 209.170 1808.100 209.695 ;
        RECT 1809.075 209.170 1809.355 210.965 ;
        RECT 1811.835 209.170 1812.115 210.965 ;
        RECT 1812.500 209.170 1812.760 209.430 ;
        RECT 1807.960 209.110 1812.760 209.170 ;
        RECT 1807.960 209.030 1812.700 209.110 ;
        RECT 1815.055 209.030 1815.460 210.965 ;
        RECT 1820.320 209.170 1820.580 209.430 ;
        RECT 1821.035 209.170 1821.315 210.965 ;
        RECT 1824.255 209.170 1824.660 210.965 ;
        RECT 1820.320 209.110 1824.660 209.170 ;
        RECT 1820.380 209.030 1824.660 209.110 ;
        RECT 1827.475 209.030 1827.880 210.965 ;
        RECT 1793.435 208.565 1793.715 209.030 ;
        RECT 1799.875 208.565 1800.155 209.030 ;
        RECT 1801.920 208.770 1802.180 209.030 ;
        RECT 1802.635 208.565 1802.915 209.030 ;
        RECT 1805.855 208.565 1806.135 209.030 ;
        RECT 1809.075 208.565 1809.355 209.030 ;
        RECT 1811.835 208.565 1812.115 209.030 ;
        RECT 1815.055 208.565 1815.335 209.030 ;
        RECT 1821.035 208.565 1821.315 209.030 ;
        RECT 1824.255 208.565 1824.535 209.030 ;
        RECT 1827.475 208.565 1827.755 209.030 ;
        RECT 1830.235 208.565 1830.515 210.965 ;
      LAYER met2 ;
        RECT 1752.085 208.285 1753.135 208.565 ;
        RECT 1753.975 208.285 1756.355 208.565 ;
        RECT 1757.195 208.285 1759.575 208.565 ;
        RECT 1760.415 208.285 1762.335 208.565 ;
        RECT 1763.175 208.285 1765.555 208.565 ;
        RECT 1766.395 208.285 1768.775 208.565 ;
        RECT 1769.615 208.285 1771.535 208.565 ;
        RECT 1772.375 208.285 1774.755 208.565 ;
        RECT 1775.595 208.285 1777.975 208.565 ;
        RECT 1778.815 208.285 1780.735 208.565 ;
        RECT 1781.575 208.285 1783.955 208.565 ;
        RECT 1784.795 208.285 1787.175 208.565 ;
        RECT 1788.015 208.285 1789.935 208.565 ;
        RECT 1790.775 208.285 1793.155 208.565 ;
        RECT 1793.995 208.285 1796.375 208.565 ;
        RECT 1797.215 208.285 1799.595 208.565 ;
        RECT 1800.435 208.285 1802.355 208.565 ;
        RECT 1803.195 208.285 1805.575 208.565 ;
        RECT 1806.415 208.285 1808.795 208.565 ;
        RECT 1809.635 208.285 1811.555 208.565 ;
        RECT 1812.395 208.285 1814.775 208.565 ;
        RECT 1815.615 208.285 1817.995 208.565 ;
        RECT 1818.835 208.285 1820.755 208.565 ;
        RECT 1821.595 208.285 1823.975 208.565 ;
        RECT 1824.815 208.285 1827.195 208.565 ;
        RECT 1828.035 208.285 1829.955 208.565 ;
        RECT 1830.795 208.285 1831.790 208.565 ;
      LAYER met2 ;
        RECT 1379.700 207.730 1380.300 207.810 ;
        RECT 1572.900 207.730 1573.500 207.810 ;
        RECT 1283.040 207.410 1283.300 207.730 ;
        RECT 1379.640 207.670 1380.360 207.730 ;
        RECT 1379.640 207.410 1379.900 207.670 ;
        RECT 1380.100 207.410 1380.360 207.670 ;
        RECT 1545.240 207.410 1545.500 207.730 ;
        RECT 1572.840 207.670 1573.560 207.730 ;
        RECT 1572.840 207.410 1573.100 207.670 ;
        RECT 1573.300 207.410 1573.560 207.670 ;
        RECT 1283.100 201.805 1283.240 207.410 ;
        RECT 1449.100 207.245 1449.360 207.390 ;
        RECT 1545.300 207.245 1545.440 207.410 ;
        RECT 1642.300 207.245 1642.560 207.390 ;
        RECT 1711.300 207.245 1711.560 207.390 ;
        RECT 1449.090 206.875 1449.370 207.245 ;
        RECT 1545.230 206.875 1545.510 207.245 ;
        RECT 1642.290 206.875 1642.570 207.245 ;
        RECT 1711.290 206.875 1711.570 207.245 ;
        RECT 1283.030 201.435 1283.310 201.805 ;
        RECT 1265.100 200.610 1265.360 200.930 ;
        RECT 1257.740 200.270 1258.000 200.590 ;
        RECT 1262.800 200.270 1263.060 200.590 ;
        RECT 1262.860 200.000 1263.000 200.270 ;
        RECT 1265.160 200.000 1265.300 200.610 ;
        RECT 667.710 174.340 691.610 200.000 ;
      LAYER met2 ;
        RECT 691.890 197.665 717.325 197.965 ;
      LAYER met2 ;
        RECT 717.605 197.945 741.505 200.000 ;
      LAYER met2 ;
        RECT 1209.085 199.080 1250.700 200.000 ;
      LAYER met2 ;
        RECT 1250.980 199.360 1251.240 200.000 ;
      LAYER met2 ;
        RECT 1251.520 199.390 1252.565 200.000 ;
      LAYER met2 ;
        RECT 1252.845 199.670 1253.495 200.000 ;
      LAYER met2 ;
        RECT 1253.775 199.390 1255.490 200.000 ;
      LAYER met2 ;
        RECT 1255.770 199.670 1256.420 200.000 ;
      LAYER met2 ;
        RECT 1256.700 199.390 1261.060 200.000 ;
        RECT 1251.520 199.080 1261.060 199.390 ;
        RECT 691.890 174.060 741.735 197.665 ;
        RECT 667.710 4.925 741.735 174.060 ;
        RECT 1209.085 196.020 1261.060 199.080 ;
        RECT 1209.085 195.735 1260.775 196.020 ;
      LAYER met2 ;
        RECT 1261.340 195.755 1261.640 200.000 ;
      LAYER met2 ;
        RECT 1261.920 198.735 1268.585 200.000 ;
      LAYER met2 ;
        RECT 1268.865 199.015 1269.445 200.000 ;
      LAYER met2 ;
        RECT 1269.725 198.735 1271.175 200.000 ;
        RECT 1261.920 198.250 1271.175 198.735 ;
        RECT 1271.995 198.250 1283.660 200.000 ;
        RECT 1261.920 196.845 1283.660 198.250 ;
        RECT 1261.920 196.485 1268.475 196.845 ;
        RECT 1273.600 196.705 1283.660 196.845 ;
        RECT 1261.920 196.215 1268.205 196.485 ;
      LAYER met2 ;
        RECT 1268.755 196.425 1273.320 196.565 ;
        RECT 1268.755 196.355 1273.650 196.425 ;
      LAYER met2 ;
        RECT 1273.930 196.375 1283.660 196.705 ;
      LAYER met2 ;
        RECT 1268.755 196.305 1273.180 196.355 ;
      LAYER met2 ;
        RECT 1261.920 196.035 1267.835 196.215 ;
      LAYER met2 ;
        RECT 1268.755 196.205 1269.115 196.305 ;
        RECT 1269.125 196.205 1269.225 196.305 ;
        RECT 1273.070 196.235 1273.305 196.305 ;
        RECT 1273.320 196.235 1273.650 196.355 ;
      LAYER met2 ;
        RECT 1262.220 195.845 1267.835 196.035 ;
      LAYER met2 ;
        RECT 1268.485 196.165 1268.755 196.205 ;
        RECT 1268.855 196.165 1269.125 196.205 ;
        RECT 1268.485 196.025 1269.125 196.165 ;
        RECT 1273.070 196.095 1273.650 196.235 ;
        RECT 1273.070 196.070 1273.305 196.095 ;
        RECT 1268.485 195.935 1268.755 196.025 ;
        RECT 1268.855 195.935 1269.125 196.025 ;
        RECT 1261.340 195.740 1261.940 195.755 ;
      LAYER met2 ;
        RECT 1209.085 195.380 1254.600 195.735 ;
      LAYER met2 ;
        RECT 1261.055 195.455 1261.940 195.740 ;
      LAYER met2 ;
        RECT 1262.220 195.735 1267.725 195.845 ;
      LAYER met2 ;
        RECT 1268.115 195.565 1268.855 195.935 ;
      LAYER met2 ;
        RECT 1269.505 195.925 1272.790 196.025 ;
        RECT 1269.405 195.790 1272.790 195.925 ;
      LAYER met2 ;
        RECT 1273.305 195.955 1273.625 196.070 ;
        RECT 1273.650 195.955 1273.995 196.095 ;
      LAYER met2 ;
        RECT 1274.275 196.030 1283.660 196.375 ;
      LAYER met2 ;
        RECT 1273.305 195.815 1273.995 195.955 ;
      LAYER met2 ;
        RECT 1269.405 195.655 1273.025 195.790 ;
      LAYER met2 ;
        RECT 1273.305 195.750 1273.625 195.815 ;
        RECT 1273.650 195.750 1273.995 195.815 ;
        RECT 1268.005 195.455 1268.485 195.565 ;
      LAYER met2 ;
        RECT 1209.085 195.050 1254.270 195.380 ;
      LAYER met2 ;
        RECT 1254.880 195.315 1268.485 195.455 ;
        RECT 1254.880 195.245 1255.235 195.315 ;
        RECT 1261.340 195.245 1261.640 195.315 ;
        RECT 1268.115 195.245 1268.485 195.315 ;
      LAYER met2 ;
        RECT 1269.135 195.470 1273.025 195.655 ;
      LAYER met2 ;
        RECT 1273.625 195.675 1273.955 195.750 ;
        RECT 1273.995 195.675 1274.265 195.750 ;
      LAYER met2 ;
        RECT 1269.135 195.285 1273.345 195.470 ;
      LAYER met2 ;
        RECT 1273.625 195.425 1274.265 195.675 ;
        RECT 1273.625 195.420 1273.955 195.425 ;
        RECT 1254.880 195.195 1268.485 195.245 ;
        RECT 1254.880 195.100 1255.235 195.195 ;
        RECT 1255.250 195.100 1255.345 195.195 ;
      LAYER met2 ;
        RECT 1268.765 195.140 1273.345 195.285 ;
      LAYER met2 ;
        RECT 1254.550 195.055 1254.880 195.100 ;
        RECT 1254.920 195.055 1255.250 195.100 ;
      LAYER met2 ;
        RECT 1209.085 189.305 1254.140 195.050 ;
      LAYER met2 ;
        RECT 1254.550 194.845 1255.250 195.055 ;
      LAYER met2 ;
        RECT 1268.765 194.915 1273.725 195.140 ;
      LAYER met2 ;
        RECT 1254.550 194.770 1254.880 194.845 ;
        RECT 1254.920 194.770 1255.250 194.845 ;
      LAYER met2 ;
        RECT 1255.625 194.820 1273.725 194.915 ;
      LAYER met2 ;
        RECT 1254.420 194.640 1254.550 194.770 ;
        RECT 1254.680 194.640 1254.920 194.770 ;
        RECT 1254.420 194.530 1254.920 194.640 ;
      LAYER met2 ;
        RECT 1209.085 189.115 1253.950 189.305 ;
        RECT 1209.085 184.635 1253.690 189.115 ;
      LAYER met2 ;
        RECT 1254.420 189.025 1254.680 194.530 ;
      LAYER met2 ;
        RECT 1255.530 194.490 1273.725 194.820 ;
        RECT 1255.200 194.250 1273.725 194.490 ;
      LAYER met2 ;
        RECT 1254.230 188.915 1254.680 189.025 ;
        RECT 1254.230 188.835 1254.420 188.915 ;
        RECT 1254.600 188.835 1254.680 188.915 ;
      LAYER met2 ;
        RECT 1254.960 191.420 1273.725 194.250 ;
        RECT 1254.960 191.080 1273.385 191.420 ;
      LAYER met2 ;
        RECT 1274.005 191.140 1274.265 195.425 ;
      LAYER met2 ;
        RECT 1254.960 190.880 1273.185 191.080 ;
      LAYER met2 ;
        RECT 1273.665 190.890 1274.265 191.140 ;
      LAYER met2 ;
        RECT 1254.960 190.550 1272.855 190.880 ;
      LAYER met2 ;
        RECT 1273.665 190.800 1274.005 190.890 ;
        RECT 1274.035 190.800 1274.265 190.890 ;
        RECT 1273.465 190.750 1273.665 190.800 ;
        RECT 1273.835 190.750 1274.035 190.800 ;
        RECT 1273.465 190.680 1274.035 190.750 ;
        RECT 1273.465 190.600 1273.665 190.680 ;
        RECT 1273.835 190.600 1274.035 190.680 ;
        RECT 1253.970 188.465 1254.600 188.835 ;
      LAYER met2 ;
        RECT 1254.960 188.555 1272.595 190.550 ;
      LAYER met2 ;
        RECT 1273.135 190.540 1273.465 190.600 ;
        RECT 1273.505 190.540 1273.835 190.600 ;
        RECT 1273.135 190.400 1273.835 190.540 ;
      LAYER met2 ;
        RECT 1274.545 190.520 1283.660 196.030 ;
      LAYER met2 ;
        RECT 1273.135 190.270 1273.465 190.400 ;
        RECT 1273.505 190.270 1273.835 190.400 ;
      LAYER met2 ;
        RECT 1274.315 190.320 1283.660 190.520 ;
        RECT 1209.085 184.300 1253.355 184.635 ;
      LAYER met2 ;
        RECT 1253.970 184.355 1254.230 188.465 ;
      LAYER met2 ;
        RECT 1254.880 188.185 1272.595 188.555 ;
        RECT 1209.085 179.225 1253.095 184.300 ;
      LAYER met2 ;
        RECT 1253.635 184.105 1254.230 184.355 ;
        RECT 1253.635 184.020 1253.970 184.105 ;
        RECT 1254.005 184.020 1254.230 184.105 ;
        RECT 1253.375 183.650 1254.005 184.020 ;
      LAYER met2 ;
        RECT 1254.510 183.740 1272.595 188.185 ;
      LAYER met2 ;
        RECT 1253.375 179.505 1253.635 183.650 ;
      LAYER met2 ;
        RECT 1254.285 183.370 1272.595 183.740 ;
        RECT 1253.915 179.225 1272.595 183.370 ;
        RECT 1209.085 172.420 1272.595 179.225 ;
      LAYER met2 ;
        RECT 1272.875 189.900 1273.505 190.270 ;
      LAYER met2 ;
        RECT 1274.115 189.990 1283.660 190.320 ;
      LAYER met2 ;
        RECT 1272.875 173.390 1273.135 189.900 ;
      LAYER met2 ;
        RECT 1273.785 189.620 1283.660 189.990 ;
        RECT 1273.415 173.670 1283.660 189.620 ;
      LAYER met2 ;
        RECT 1272.875 172.700 1273.350 173.390 ;
      LAYER met2 ;
        RECT 1209.085 172.345 1272.810 172.420 ;
        RECT 1209.085 169.195 1272.595 172.345 ;
      LAYER met2 ;
        RECT 1273.090 172.065 1273.350 172.700 ;
        RECT 1272.875 171.855 1273.350 172.065 ;
        RECT 1272.875 171.850 1273.090 171.855 ;
        RECT 1272.875 171.375 1273.350 171.850 ;
      LAYER met2 ;
        RECT 1209.085 169.050 1272.450 169.195 ;
        RECT 1209.085 168.825 1272.225 169.050 ;
      LAYER met2 ;
        RECT 1272.875 168.915 1273.135 171.375 ;
      LAYER met2 ;
        RECT 1273.630 171.095 1283.660 173.670 ;
        RECT 1209.085 164.260 1272.200 168.825 ;
      LAYER met2 ;
        RECT 1272.730 168.770 1273.135 168.915 ;
        RECT 1272.505 168.735 1272.730 168.770 ;
        RECT 1272.875 168.735 1273.135 168.770 ;
        RECT 1272.505 168.665 1273.135 168.735 ;
        RECT 1272.505 168.545 1272.730 168.665 ;
        RECT 1272.875 168.545 1273.135 168.665 ;
        RECT 1272.480 168.520 1272.505 168.545 ;
        RECT 1272.740 168.520 1272.875 168.545 ;
        RECT 1272.480 168.410 1272.875 168.520 ;
      LAYER met2 ;
        RECT 1209.085 163.440 1271.570 164.260 ;
      LAYER met2 ;
        RECT 1272.480 163.980 1272.740 168.410 ;
      LAYER met2 ;
        RECT 1273.415 168.265 1283.660 171.095 ;
        RECT 1273.155 168.130 1283.660 168.265 ;
      LAYER met2 ;
        RECT 1271.850 163.720 1272.740 163.980 ;
      LAYER met2 ;
        RECT 1273.020 163.440 1283.660 168.130 ;
        RECT 1209.085 0.790 1283.660 163.440 ;
        RECT 1752.085 0.000 1831.790 208.285 ;
      LAYER met2 ;
        RECT 2304.760 200.445 2304.900 221.690 ;
        RECT 2348.920 221.670 2349.060 228.150 ;
        RECT 2370.480 227.810 2370.740 228.130 ;
        RECT 2325.400 221.350 2325.660 221.670 ;
        RECT 2348.860 221.350 2349.120 221.670 ;
        RECT 2304.690 200.075 2304.970 200.445 ;
        RECT 2304.760 198.550 2304.900 200.075 ;
        RECT 2325.460 199.765 2325.600 221.350 ;
        RECT 2370.540 221.330 2370.680 227.810 ;
        RECT 2353.460 221.010 2353.720 221.330 ;
        RECT 2370.480 221.010 2370.740 221.330 ;
        RECT 2332.300 220.670 2332.560 220.990 ;
        RECT 2325.390 199.395 2325.670 199.765 ;
        RECT 2299.180 198.230 2299.440 198.550 ;
        RECT 2304.700 198.230 2304.960 198.550 ;
        RECT 2299.240 198.000 2299.380 198.230 ;
        RECT 2332.360 198.000 2332.500 220.670 ;
        RECT 2345.630 213.675 2345.910 214.045 ;
        RECT 2337.810 200.075 2338.090 200.445 ;
        RECT 2337.880 199.085 2338.020 200.075 ;
        RECT 2345.700 199.085 2345.840 213.675 ;
        RECT 2337.810 198.715 2338.090 199.085 ;
        RECT 2345.630 198.715 2345.910 199.085 ;
        RECT 2353.520 198.000 2353.660 221.010 ;
        RECT 2911.960 220.990 2912.100 228.490 ;
        RECT 3367.360 228.470 3367.500 741.210 ;
        RECT 3367.300 228.150 3367.560 228.470 ;
        RECT 3368.280 228.130 3368.420 788.470 ;
        RECT 3368.740 741.530 3368.880 896.930 ;
        RECT 3368.680 741.210 3368.940 741.530 ;
        RECT 3373.800 228.810 3373.940 4374.450 ;
        RECT 3390.360 4364.085 3390.500 4380.300 ;
        RECT 3390.290 4363.715 3390.570 4364.085 ;
      LAYER met2 ;
        RECT 3379.435 3849.795 3588.000 3850.790 ;
      LAYER met2 ;
        RECT 3377.035 3849.235 3379.435 3849.515 ;
      LAYER met2 ;
        RECT 3379.715 3848.955 3588.000 3849.795 ;
        RECT 3379.435 3847.035 3588.000 3848.955 ;
        RECT 3379.715 3846.195 3588.000 3847.035 ;
        RECT 3379.435 3843.815 3588.000 3846.195 ;
        RECT 3379.715 3842.975 3588.000 3843.815 ;
        RECT 3379.435 3840.595 3588.000 3842.975 ;
        RECT 3379.715 3839.755 3588.000 3840.595 ;
        RECT 3379.435 3837.835 3588.000 3839.755 ;
        RECT 3379.715 3836.995 3588.000 3837.835 ;
      LAYER met2 ;
        RECT 3376.960 3836.570 3377.220 3836.890 ;
        RECT 3377.020 3834.335 3377.160 3836.570 ;
      LAYER met2 ;
        RECT 3379.435 3834.615 3588.000 3836.995 ;
      LAYER met2 ;
        RECT 3377.020 3834.180 3379.435 3834.335 ;
        RECT 3377.035 3834.055 3379.435 3834.180 ;
      LAYER met2 ;
        RECT 3379.715 3833.775 3588.000 3834.615 ;
        RECT 3379.435 3831.395 3588.000 3833.775 ;
        RECT 3379.715 3830.555 3588.000 3831.395 ;
        RECT 3379.435 3828.635 3588.000 3830.555 ;
        RECT 3379.715 3827.795 3588.000 3828.635 ;
        RECT 3379.435 3825.415 3588.000 3827.795 ;
        RECT 3379.715 3824.575 3588.000 3825.415 ;
        RECT 3379.435 3822.195 3588.000 3824.575 ;
        RECT 3379.715 3821.355 3588.000 3822.195 ;
        RECT 3379.435 3819.435 3588.000 3821.355 ;
        RECT 3379.715 3818.595 3588.000 3819.435 ;
        RECT 3379.435 3816.215 3588.000 3818.595 ;
        RECT 3379.715 3815.375 3588.000 3816.215 ;
        RECT 3379.435 3812.995 3588.000 3815.375 ;
      LAYER met2 ;
        RECT 3377.035 3812.645 3379.435 3812.715 ;
        RECT 3376.560 3812.505 3379.435 3812.645 ;
        RECT 3376.560 3772.625 3376.700 3812.505 ;
        RECT 3377.035 3812.435 3379.435 3812.505 ;
      LAYER met2 ;
        RECT 3379.715 3812.155 3588.000 3812.995 ;
        RECT 3379.435 3809.775 3588.000 3812.155 ;
        RECT 3379.715 3808.935 3588.000 3809.775 ;
        RECT 3379.435 3807.015 3588.000 3808.935 ;
        RECT 3379.715 3806.175 3588.000 3807.015 ;
        RECT 3379.435 3803.795 3588.000 3806.175 ;
        RECT 3379.715 3802.955 3588.000 3803.795 ;
        RECT 3379.435 3800.575 3588.000 3802.955 ;
        RECT 3379.715 3799.735 3588.000 3800.575 ;
        RECT 3379.435 3797.815 3588.000 3799.735 ;
      LAYER met2 ;
        RECT 3377.035 3797.255 3379.435 3797.535 ;
      LAYER met2 ;
        RECT 3379.715 3796.975 3588.000 3797.815 ;
        RECT 3379.435 3794.595 3588.000 3796.975 ;
        RECT 3379.715 3793.755 3588.000 3794.595 ;
        RECT 3379.435 3791.375 3588.000 3793.755 ;
      LAYER met2 ;
        RECT 3377.035 3790.815 3379.435 3791.095 ;
      LAYER met2 ;
        RECT 3379.715 3790.535 3588.000 3791.375 ;
        RECT 3379.435 3788.615 3588.000 3790.535 ;
      LAYER met2 ;
        RECT 3377.035 3788.055 3379.435 3788.335 ;
      LAYER met2 ;
        RECT 3379.715 3787.775 3588.000 3788.615 ;
        RECT 3379.435 3785.395 3588.000 3787.775 ;
        RECT 3379.715 3784.555 3588.000 3785.395 ;
        RECT 3379.435 3782.175 3588.000 3784.555 ;
      LAYER met2 ;
        RECT 3377.035 3781.820 3379.435 3781.895 ;
        RECT 3377.020 3781.615 3379.435 3781.820 ;
        RECT 3377.020 3779.770 3377.160 3781.615 ;
      LAYER met2 ;
        RECT 3379.715 3781.335 3588.000 3782.175 ;
      LAYER met2 ;
        RECT 3376.960 3779.450 3377.220 3779.770 ;
      LAYER met2 ;
        RECT 3379.435 3779.415 3588.000 3781.335 ;
      LAYER met2 ;
        RECT 3377.035 3778.855 3379.435 3779.135 ;
      LAYER met2 ;
        RECT 3379.715 3778.575 3588.000 3779.415 ;
        RECT 3379.435 3776.195 3588.000 3778.575 ;
        RECT 3379.715 3775.355 3588.000 3776.195 ;
        RECT 3379.435 3772.975 3588.000 3775.355 ;
      LAYER met2 ;
        RECT 3377.035 3772.625 3379.435 3772.695 ;
        RECT 3376.560 3772.485 3379.435 3772.625 ;
        RECT 3377.035 3772.415 3379.435 3772.485 ;
      LAYER met2 ;
        RECT 3379.715 3772.135 3588.000 3772.975 ;
        RECT 3379.435 3771.085 3588.000 3772.135 ;
        RECT 3379.435 3241.795 3588.000 3242.790 ;
      LAYER met2 ;
        RECT 3377.035 3241.235 3379.435 3241.515 ;
      LAYER met2 ;
        RECT 3379.715 3240.955 3588.000 3241.795 ;
        RECT 3379.435 3239.035 3588.000 3240.955 ;
        RECT 3379.715 3238.195 3588.000 3239.035 ;
        RECT 3379.435 3235.815 3588.000 3238.195 ;
        RECT 3379.715 3234.975 3588.000 3235.815 ;
        RECT 3379.435 3232.595 3588.000 3234.975 ;
        RECT 3379.715 3231.755 3588.000 3232.595 ;
        RECT 3379.435 3229.835 3588.000 3231.755 ;
        RECT 3379.715 3228.995 3588.000 3229.835 ;
      LAYER met2 ;
        RECT 3376.960 3228.650 3377.220 3228.970 ;
        RECT 3377.020 3226.335 3377.160 3228.650 ;
      LAYER met2 ;
        RECT 3379.435 3226.615 3588.000 3228.995 ;
      LAYER met2 ;
        RECT 3377.020 3226.260 3379.435 3226.335 ;
        RECT 3377.035 3226.055 3379.435 3226.260 ;
      LAYER met2 ;
        RECT 3379.715 3225.775 3588.000 3226.615 ;
        RECT 3379.435 3223.395 3588.000 3225.775 ;
        RECT 3379.715 3222.555 3588.000 3223.395 ;
        RECT 3379.435 3220.635 3588.000 3222.555 ;
        RECT 3379.715 3219.795 3588.000 3220.635 ;
        RECT 3379.435 3217.415 3588.000 3219.795 ;
        RECT 3379.715 3216.575 3588.000 3217.415 ;
        RECT 3379.435 3214.195 3588.000 3216.575 ;
        RECT 3379.715 3213.355 3588.000 3214.195 ;
        RECT 3379.435 3211.435 3588.000 3213.355 ;
        RECT 3379.715 3210.595 3588.000 3211.435 ;
        RECT 3379.435 3208.215 3588.000 3210.595 ;
        RECT 3379.715 3207.375 3588.000 3208.215 ;
        RECT 3379.435 3204.995 3588.000 3207.375 ;
      LAYER met2 ;
        RECT 3377.035 3204.570 3379.435 3204.715 ;
        RECT 3376.560 3204.435 3379.435 3204.570 ;
        RECT 3376.560 3204.430 3377.090 3204.435 ;
        RECT 3376.560 3164.625 3376.700 3204.430 ;
      LAYER met2 ;
        RECT 3379.715 3204.155 3588.000 3204.995 ;
        RECT 3379.435 3201.775 3588.000 3204.155 ;
        RECT 3379.715 3200.935 3588.000 3201.775 ;
        RECT 3379.435 3199.015 3588.000 3200.935 ;
        RECT 3379.715 3198.175 3588.000 3199.015 ;
        RECT 3379.435 3195.795 3588.000 3198.175 ;
        RECT 3379.715 3194.955 3588.000 3195.795 ;
        RECT 3379.435 3192.575 3588.000 3194.955 ;
        RECT 3379.715 3191.735 3588.000 3192.575 ;
        RECT 3379.435 3189.815 3588.000 3191.735 ;
      LAYER met2 ;
        RECT 3377.035 3189.255 3379.435 3189.535 ;
      LAYER met2 ;
        RECT 3379.715 3188.975 3588.000 3189.815 ;
        RECT 3379.435 3186.595 3588.000 3188.975 ;
        RECT 3379.715 3185.755 3588.000 3186.595 ;
        RECT 3379.435 3183.375 3588.000 3185.755 ;
      LAYER met2 ;
        RECT 3377.035 3182.815 3379.435 3183.095 ;
      LAYER met2 ;
        RECT 3379.715 3182.535 3588.000 3183.375 ;
        RECT 3379.435 3180.615 3588.000 3182.535 ;
      LAYER met2 ;
        RECT 3377.035 3180.055 3379.435 3180.335 ;
      LAYER met2 ;
        RECT 3379.715 3179.775 3588.000 3180.615 ;
        RECT 3379.435 3177.395 3588.000 3179.775 ;
        RECT 3379.715 3176.555 3588.000 3177.395 ;
        RECT 3379.435 3174.175 3588.000 3176.555 ;
      LAYER met2 ;
        RECT 3377.035 3173.755 3379.435 3173.895 ;
        RECT 3377.020 3173.615 3379.435 3173.755 ;
        RECT 3377.020 3171.850 3377.160 3173.615 ;
      LAYER met2 ;
        RECT 3379.715 3173.335 3588.000 3174.175 ;
      LAYER met2 ;
        RECT 3376.960 3171.530 3377.220 3171.850 ;
      LAYER met2 ;
        RECT 3379.435 3171.415 3588.000 3173.335 ;
      LAYER met2 ;
        RECT 3377.035 3170.855 3379.435 3171.135 ;
      LAYER met2 ;
        RECT 3379.715 3170.575 3588.000 3171.415 ;
        RECT 3379.435 3168.195 3588.000 3170.575 ;
        RECT 3379.715 3167.355 3588.000 3168.195 ;
        RECT 3379.435 3164.975 3588.000 3167.355 ;
      LAYER met2 ;
        RECT 3377.035 3164.625 3379.435 3164.695 ;
        RECT 3376.560 3164.485 3379.435 3164.625 ;
        RECT 3377.035 3164.415 3379.435 3164.485 ;
      LAYER met2 ;
        RECT 3379.715 3164.135 3588.000 3164.975 ;
        RECT 3379.435 3163.085 3588.000 3164.135 ;
        RECT 3379.435 2632.795 3588.000 2633.790 ;
      LAYER met2 ;
        RECT 3377.035 2632.235 3379.435 2632.515 ;
      LAYER met2 ;
        RECT 3379.715 2631.955 3588.000 2632.795 ;
        RECT 3379.435 2630.035 3588.000 2631.955 ;
        RECT 3379.715 2629.195 3588.000 2630.035 ;
        RECT 3379.435 2626.815 3588.000 2629.195 ;
        RECT 3379.715 2625.975 3588.000 2626.815 ;
        RECT 3379.435 2623.595 3588.000 2625.975 ;
        RECT 3379.715 2622.755 3588.000 2623.595 ;
        RECT 3379.435 2620.835 3588.000 2622.755 ;
        RECT 3379.715 2619.995 3588.000 2620.835 ;
        RECT 3379.435 2617.615 3588.000 2619.995 ;
      LAYER met2 ;
        RECT 3377.035 2617.195 3379.435 2617.335 ;
        RECT 3377.020 2617.055 3379.435 2617.195 ;
        RECT 3377.020 2614.590 3377.160 2617.055 ;
      LAYER met2 ;
        RECT 3379.715 2616.775 3588.000 2617.615 ;
      LAYER met2 ;
        RECT 3376.960 2614.270 3377.220 2614.590 ;
      LAYER met2 ;
        RECT 3379.435 2614.395 3588.000 2616.775 ;
        RECT 3379.715 2613.555 3588.000 2614.395 ;
        RECT 3379.435 2611.635 3588.000 2613.555 ;
        RECT 3379.715 2610.795 3588.000 2611.635 ;
        RECT 3379.435 2608.415 3588.000 2610.795 ;
        RECT 3379.715 2607.575 3588.000 2608.415 ;
        RECT 3379.435 2605.195 3588.000 2607.575 ;
        RECT 3379.715 2604.355 3588.000 2605.195 ;
        RECT 3379.435 2602.435 3588.000 2604.355 ;
        RECT 3379.715 2601.595 3588.000 2602.435 ;
        RECT 3379.435 2599.215 3588.000 2601.595 ;
        RECT 3379.715 2598.375 3588.000 2599.215 ;
        RECT 3379.435 2595.995 3588.000 2598.375 ;
      LAYER met2 ;
        RECT 3377.035 2595.645 3379.435 2595.715 ;
        RECT 3376.560 2595.505 3379.435 2595.645 ;
        RECT 3376.560 2555.625 3376.700 2595.505 ;
        RECT 3377.035 2595.435 3379.435 2595.505 ;
      LAYER met2 ;
        RECT 3379.715 2595.155 3588.000 2595.995 ;
        RECT 3379.435 2592.775 3588.000 2595.155 ;
        RECT 3379.715 2591.935 3588.000 2592.775 ;
        RECT 3379.435 2590.015 3588.000 2591.935 ;
        RECT 3379.715 2589.175 3588.000 2590.015 ;
        RECT 3379.435 2586.795 3588.000 2589.175 ;
        RECT 3379.715 2585.955 3588.000 2586.795 ;
        RECT 3379.435 2583.575 3588.000 2585.955 ;
        RECT 3379.715 2582.735 3588.000 2583.575 ;
        RECT 3379.435 2580.815 3588.000 2582.735 ;
      LAYER met2 ;
        RECT 3377.035 2580.255 3379.435 2580.535 ;
      LAYER met2 ;
        RECT 3379.715 2579.975 3588.000 2580.815 ;
        RECT 3379.435 2577.595 3588.000 2579.975 ;
        RECT 3379.715 2576.755 3588.000 2577.595 ;
        RECT 3379.435 2574.375 3588.000 2576.755 ;
      LAYER met2 ;
        RECT 3377.035 2573.815 3379.435 2574.095 ;
      LAYER met2 ;
        RECT 3379.715 2573.535 3588.000 2574.375 ;
        RECT 3379.435 2571.615 3588.000 2573.535 ;
      LAYER met2 ;
        RECT 3377.035 2571.055 3379.435 2571.335 ;
      LAYER met2 ;
        RECT 3379.715 2570.775 3588.000 2571.615 ;
        RECT 3379.435 2568.395 3588.000 2570.775 ;
        RECT 3379.715 2567.555 3588.000 2568.395 ;
      LAYER met2 ;
        RECT 3376.960 2565.310 3377.220 2565.630 ;
        RECT 3377.020 2564.895 3377.160 2565.310 ;
      LAYER met2 ;
        RECT 3379.435 2565.175 3588.000 2567.555 ;
      LAYER met2 ;
        RECT 3377.020 2564.620 3379.435 2564.895 ;
        RECT 3377.035 2564.615 3379.435 2564.620 ;
      LAYER met2 ;
        RECT 3379.715 2564.335 3588.000 2565.175 ;
        RECT 3379.435 2562.415 3588.000 2564.335 ;
      LAYER met2 ;
        RECT 3377.035 2561.855 3379.435 2562.135 ;
      LAYER met2 ;
        RECT 3379.715 2561.575 3588.000 2562.415 ;
        RECT 3379.435 2559.195 3588.000 2561.575 ;
        RECT 3379.715 2558.355 3588.000 2559.195 ;
        RECT 3379.435 2555.975 3588.000 2558.355 ;
      LAYER met2 ;
        RECT 3377.035 2555.625 3379.435 2555.695 ;
        RECT 3376.560 2555.485 3379.435 2555.625 ;
        RECT 3377.035 2555.415 3379.435 2555.485 ;
      LAYER met2 ;
        RECT 3379.715 2555.135 3588.000 2555.975 ;
        RECT 3379.435 2554.085 3588.000 2555.135 ;
        RECT 3379.435 2023.795 3588.000 2024.790 ;
      LAYER met2 ;
        RECT 3377.035 2023.235 3379.435 2023.515 ;
      LAYER met2 ;
        RECT 3379.715 2022.955 3588.000 2023.795 ;
        RECT 3379.435 2021.035 3588.000 2022.955 ;
        RECT 3379.715 2020.195 3588.000 2021.035 ;
        RECT 3379.435 2017.815 3588.000 2020.195 ;
        RECT 3379.715 2016.975 3588.000 2017.815 ;
        RECT 3379.435 2014.595 3588.000 2016.975 ;
        RECT 3379.715 2013.755 3588.000 2014.595 ;
        RECT 3379.435 2011.835 3588.000 2013.755 ;
        RECT 3379.715 2010.995 3588.000 2011.835 ;
        RECT 3379.435 2008.615 3588.000 2010.995 ;
      LAYER met2 ;
        RECT 3377.035 2008.195 3379.435 2008.335 ;
        RECT 3377.020 2008.055 3379.435 2008.195 ;
        RECT 3377.020 2007.010 3377.160 2008.055 ;
      LAYER met2 ;
        RECT 3379.715 2007.775 3588.000 2008.615 ;
      LAYER met2 ;
        RECT 3376.960 2006.690 3377.220 2007.010 ;
      LAYER met2 ;
        RECT 3379.435 2005.395 3588.000 2007.775 ;
        RECT 3379.715 2004.555 3588.000 2005.395 ;
        RECT 3379.435 2002.635 3588.000 2004.555 ;
        RECT 3379.715 2001.795 3588.000 2002.635 ;
        RECT 3379.435 1999.415 3588.000 2001.795 ;
        RECT 3379.715 1998.575 3588.000 1999.415 ;
        RECT 3379.435 1996.195 3588.000 1998.575 ;
        RECT 3379.715 1995.355 3588.000 1996.195 ;
        RECT 3379.435 1993.435 3588.000 1995.355 ;
        RECT 3379.715 1992.595 3588.000 1993.435 ;
        RECT 3379.435 1990.215 3588.000 1992.595 ;
        RECT 3379.715 1989.375 3588.000 1990.215 ;
        RECT 3379.435 1986.995 3588.000 1989.375 ;
      LAYER met2 ;
        RECT 3377.035 1986.690 3379.435 1986.715 ;
        RECT 3376.560 1986.550 3379.435 1986.690 ;
        RECT 3376.560 1946.570 3376.700 1986.550 ;
        RECT 3377.035 1986.435 3379.435 1986.550 ;
      LAYER met2 ;
        RECT 3379.715 1986.155 3588.000 1986.995 ;
        RECT 3379.435 1983.775 3588.000 1986.155 ;
        RECT 3379.715 1982.935 3588.000 1983.775 ;
        RECT 3379.435 1981.015 3588.000 1982.935 ;
        RECT 3379.715 1980.175 3588.000 1981.015 ;
        RECT 3379.435 1977.795 3588.000 1980.175 ;
        RECT 3379.715 1976.955 3588.000 1977.795 ;
        RECT 3379.435 1974.575 3588.000 1976.955 ;
        RECT 3379.715 1973.735 3588.000 1974.575 ;
        RECT 3379.435 1971.815 3588.000 1973.735 ;
      LAYER met2 ;
        RECT 3377.035 1971.255 3379.435 1971.535 ;
      LAYER met2 ;
        RECT 3379.715 1970.975 3588.000 1971.815 ;
        RECT 3379.435 1968.595 3588.000 1970.975 ;
        RECT 3379.715 1967.755 3588.000 1968.595 ;
        RECT 3379.435 1965.375 3588.000 1967.755 ;
      LAYER met2 ;
        RECT 3377.035 1964.815 3379.435 1965.095 ;
      LAYER met2 ;
        RECT 3379.715 1964.535 3588.000 1965.375 ;
        RECT 3379.435 1962.615 3588.000 1964.535 ;
      LAYER met2 ;
        RECT 3377.035 1962.055 3379.435 1962.335 ;
      LAYER met2 ;
        RECT 3379.715 1961.775 3588.000 1962.615 ;
        RECT 3379.435 1959.395 3588.000 1961.775 ;
        RECT 3379.715 1958.555 3588.000 1959.395 ;
      LAYER met2 ;
        RECT 3376.960 1958.070 3377.220 1958.390 ;
        RECT 3377.020 1955.895 3377.160 1958.070 ;
      LAYER met2 ;
        RECT 3379.435 1956.175 3588.000 1958.555 ;
      LAYER met2 ;
        RECT 3377.020 1955.755 3379.435 1955.895 ;
        RECT 3377.035 1955.615 3379.435 1955.755 ;
      LAYER met2 ;
        RECT 3379.715 1955.335 3588.000 1956.175 ;
        RECT 3379.435 1953.415 3588.000 1955.335 ;
      LAYER met2 ;
        RECT 3377.035 1952.855 3379.435 1953.135 ;
      LAYER met2 ;
        RECT 3379.715 1952.575 3588.000 1953.415 ;
        RECT 3379.435 1950.195 3588.000 1952.575 ;
        RECT 3379.715 1949.355 3588.000 1950.195 ;
        RECT 3379.435 1946.975 3588.000 1949.355 ;
      LAYER met2 ;
        RECT 3377.035 1946.570 3379.435 1946.695 ;
        RECT 3376.560 1946.430 3379.435 1946.570 ;
        RECT 3377.035 1946.415 3379.435 1946.430 ;
      LAYER met2 ;
        RECT 3379.715 1946.135 3588.000 1946.975 ;
        RECT 3379.435 1945.085 3588.000 1946.135 ;
      LAYER met2 ;
        RECT 3376.500 1418.830 3376.760 1419.150 ;
        RECT 3376.560 1402.570 3376.700 1418.830 ;
      LAYER met2 ;
        RECT 3379.435 1415.795 3588.000 1416.790 ;
      LAYER met2 ;
        RECT 3377.035 1415.235 3379.435 1415.515 ;
      LAYER met2 ;
        RECT 3379.715 1414.955 3588.000 1415.795 ;
        RECT 3379.435 1413.035 3588.000 1414.955 ;
        RECT 3379.715 1412.195 3588.000 1413.035 ;
        RECT 3379.435 1409.815 3588.000 1412.195 ;
        RECT 3379.715 1408.975 3588.000 1409.815 ;
        RECT 3379.435 1406.595 3588.000 1408.975 ;
        RECT 3379.715 1405.755 3588.000 1406.595 ;
        RECT 3379.435 1403.835 3588.000 1405.755 ;
        RECT 3379.715 1402.995 3588.000 1403.835 ;
      LAYER met2 ;
        RECT 3376.560 1402.430 3377.160 1402.570 ;
        RECT 3377.020 1400.335 3377.160 1402.430 ;
      LAYER met2 ;
        RECT 3379.435 1400.615 3588.000 1402.995 ;
      LAYER met2 ;
        RECT 3377.020 1400.195 3379.435 1400.335 ;
        RECT 3377.035 1400.055 3379.435 1400.195 ;
      LAYER met2 ;
        RECT 3379.715 1399.775 3588.000 1400.615 ;
        RECT 3379.435 1397.395 3588.000 1399.775 ;
        RECT 3379.715 1396.555 3588.000 1397.395 ;
        RECT 3379.435 1394.635 3588.000 1396.555 ;
        RECT 3379.715 1393.795 3588.000 1394.635 ;
        RECT 3379.435 1391.415 3588.000 1393.795 ;
        RECT 3379.715 1390.575 3588.000 1391.415 ;
        RECT 3379.435 1388.195 3588.000 1390.575 ;
        RECT 3379.715 1387.355 3588.000 1388.195 ;
        RECT 3379.435 1385.435 3588.000 1387.355 ;
        RECT 3379.715 1384.595 3588.000 1385.435 ;
        RECT 3379.435 1382.215 3588.000 1384.595 ;
        RECT 3379.715 1381.375 3588.000 1382.215 ;
        RECT 3379.435 1378.995 3588.000 1381.375 ;
      LAYER met2 ;
        RECT 3377.035 1378.700 3379.435 1378.715 ;
        RECT 3377.020 1378.435 3379.435 1378.700 ;
        RECT 3377.020 1376.050 3377.160 1378.435 ;
      LAYER met2 ;
        RECT 3379.715 1378.155 3588.000 1378.995 ;
      LAYER met2 ;
        RECT 3376.560 1375.910 3377.160 1376.050 ;
        RECT 3376.560 1338.650 3376.700 1375.910 ;
      LAYER met2 ;
        RECT 3379.435 1375.775 3588.000 1378.155 ;
        RECT 3379.715 1374.935 3588.000 1375.775 ;
        RECT 3379.435 1373.015 3588.000 1374.935 ;
        RECT 3379.715 1372.175 3588.000 1373.015 ;
        RECT 3379.435 1369.795 3588.000 1372.175 ;
        RECT 3379.715 1368.955 3588.000 1369.795 ;
        RECT 3379.435 1366.575 3588.000 1368.955 ;
        RECT 3379.715 1365.735 3588.000 1366.575 ;
        RECT 3379.435 1363.815 3588.000 1365.735 ;
      LAYER met2 ;
        RECT 3377.035 1363.255 3379.435 1363.535 ;
      LAYER met2 ;
        RECT 3379.715 1362.975 3588.000 1363.815 ;
        RECT 3379.435 1360.595 3588.000 1362.975 ;
        RECT 3379.715 1359.755 3588.000 1360.595 ;
        RECT 3379.435 1357.375 3588.000 1359.755 ;
      LAYER met2 ;
        RECT 3377.035 1356.815 3379.435 1357.095 ;
      LAYER met2 ;
        RECT 3379.715 1356.535 3588.000 1357.375 ;
        RECT 3379.435 1354.615 3588.000 1356.535 ;
      LAYER met2 ;
        RECT 3377.035 1354.055 3379.435 1354.335 ;
      LAYER met2 ;
        RECT 3379.715 1353.775 3588.000 1354.615 ;
        RECT 3379.435 1351.395 3588.000 1353.775 ;
        RECT 3379.715 1350.555 3588.000 1351.395 ;
        RECT 3379.435 1348.175 3588.000 1350.555 ;
      LAYER met2 ;
        RECT 3377.035 1347.755 3379.435 1347.895 ;
        RECT 3377.020 1347.615 3379.435 1347.755 ;
        RECT 3377.020 1345.710 3377.160 1347.615 ;
      LAYER met2 ;
        RECT 3379.715 1347.335 3588.000 1348.175 ;
      LAYER met2 ;
        RECT 3376.960 1345.390 3377.220 1345.710 ;
      LAYER met2 ;
        RECT 3379.435 1345.415 3588.000 1347.335 ;
      LAYER met2 ;
        RECT 3377.035 1344.855 3379.435 1345.135 ;
      LAYER met2 ;
        RECT 3379.715 1344.575 3588.000 1345.415 ;
        RECT 3379.435 1342.195 3588.000 1344.575 ;
        RECT 3379.715 1341.355 3588.000 1342.195 ;
        RECT 3379.435 1338.975 3588.000 1341.355 ;
      LAYER met2 ;
        RECT 3377.035 1338.650 3379.435 1338.695 ;
        RECT 3376.560 1338.510 3379.435 1338.650 ;
        RECT 3377.035 1338.415 3379.435 1338.510 ;
      LAYER met2 ;
        RECT 3379.715 1338.135 3588.000 1338.975 ;
        RECT 3379.435 1337.085 3588.000 1338.135 ;
        RECT 3379.435 806.795 3588.000 807.790 ;
      LAYER met2 ;
        RECT 3377.035 806.235 3379.435 806.515 ;
      LAYER met2 ;
        RECT 3379.715 805.955 3588.000 806.795 ;
        RECT 3379.435 804.035 3588.000 805.955 ;
        RECT 3379.715 803.195 3588.000 804.035 ;
        RECT 3379.435 800.815 3588.000 803.195 ;
        RECT 3379.715 799.975 3588.000 800.815 ;
        RECT 3379.435 797.595 3588.000 799.975 ;
        RECT 3379.715 796.755 3588.000 797.595 ;
        RECT 3379.435 794.835 3588.000 796.755 ;
        RECT 3379.715 793.995 3588.000 794.835 ;
        RECT 3379.435 791.615 3588.000 793.995 ;
      LAYER met2 ;
        RECT 3377.035 791.180 3379.435 791.335 ;
        RECT 3377.020 791.055 3379.435 791.180 ;
        RECT 3377.020 788.790 3377.160 791.055 ;
      LAYER met2 ;
        RECT 3379.715 790.775 3588.000 791.615 ;
      LAYER met2 ;
        RECT 3376.960 788.470 3377.220 788.790 ;
      LAYER met2 ;
        RECT 3379.435 788.395 3588.000 790.775 ;
        RECT 3379.715 787.555 3588.000 788.395 ;
        RECT 3379.435 785.635 3588.000 787.555 ;
        RECT 3379.715 784.795 3588.000 785.635 ;
        RECT 3379.435 782.415 3588.000 784.795 ;
        RECT 3379.715 781.575 3588.000 782.415 ;
        RECT 3379.435 779.195 3588.000 781.575 ;
        RECT 3379.715 778.355 3588.000 779.195 ;
        RECT 3379.435 776.435 3588.000 778.355 ;
        RECT 3379.715 775.595 3588.000 776.435 ;
        RECT 3379.435 773.215 3588.000 775.595 ;
        RECT 3379.715 772.375 3588.000 773.215 ;
        RECT 3379.435 769.995 3588.000 772.375 ;
      LAYER met2 ;
        RECT 3377.035 769.645 3379.435 769.715 ;
        RECT 3376.560 769.505 3379.435 769.645 ;
        RECT 3376.560 729.625 3376.700 769.505 ;
        RECT 3377.035 769.435 3379.435 769.505 ;
      LAYER met2 ;
        RECT 3379.715 769.155 3588.000 769.995 ;
        RECT 3379.435 766.775 3588.000 769.155 ;
        RECT 3379.715 765.935 3588.000 766.775 ;
        RECT 3379.435 764.015 3588.000 765.935 ;
        RECT 3379.715 763.175 3588.000 764.015 ;
        RECT 3379.435 760.795 3588.000 763.175 ;
        RECT 3379.715 759.955 3588.000 760.795 ;
        RECT 3379.435 757.575 3588.000 759.955 ;
        RECT 3379.715 756.735 3588.000 757.575 ;
        RECT 3379.435 754.815 3588.000 756.735 ;
      LAYER met2 ;
        RECT 3377.035 754.255 3379.435 754.535 ;
      LAYER met2 ;
        RECT 3379.715 753.975 3588.000 754.815 ;
        RECT 3379.435 751.595 3588.000 753.975 ;
        RECT 3379.715 750.755 3588.000 751.595 ;
        RECT 3379.435 748.375 3588.000 750.755 ;
      LAYER met2 ;
        RECT 3377.035 747.815 3379.435 748.095 ;
      LAYER met2 ;
        RECT 3379.715 747.535 3588.000 748.375 ;
        RECT 3379.435 745.615 3588.000 747.535 ;
      LAYER met2 ;
        RECT 3377.035 745.055 3379.435 745.335 ;
      LAYER met2 ;
        RECT 3379.715 744.775 3588.000 745.615 ;
        RECT 3379.435 742.395 3588.000 744.775 ;
        RECT 3379.715 741.555 3588.000 742.395 ;
      LAYER met2 ;
        RECT 3376.960 741.210 3377.220 741.530 ;
        RECT 3377.020 738.895 3377.160 741.210 ;
      LAYER met2 ;
        RECT 3379.435 739.175 3588.000 741.555 ;
      LAYER met2 ;
        RECT 3377.020 738.820 3379.435 738.895 ;
        RECT 3377.035 738.615 3379.435 738.820 ;
      LAYER met2 ;
        RECT 3379.715 738.335 3588.000 739.175 ;
        RECT 3379.435 736.415 3588.000 738.335 ;
      LAYER met2 ;
        RECT 3377.035 735.855 3379.435 736.135 ;
      LAYER met2 ;
        RECT 3379.715 735.575 3588.000 736.415 ;
        RECT 3379.435 733.195 3588.000 735.575 ;
        RECT 3379.715 732.355 3588.000 733.195 ;
        RECT 3379.435 729.975 3588.000 732.355 ;
      LAYER met2 ;
        RECT 3377.035 729.625 3379.435 729.695 ;
        RECT 3376.560 729.485 3379.435 729.625 ;
        RECT 3377.035 729.415 3379.435 729.485 ;
      LAYER met2 ;
        RECT 3379.715 729.135 3588.000 729.975 ;
        RECT 3379.435 728.085 3588.000 729.135 ;
      LAYER met2 ;
        RECT 3384.310 482.275 3384.590 482.645 ;
        RECT 3384.380 386.765 3384.520 482.275 ;
        RECT 3384.310 386.395 3384.590 386.765 ;
        RECT 3383.390 385.715 3383.670 386.085 ;
        RECT 3383.460 290.205 3383.600 385.715 ;
        RECT 3383.390 289.835 3383.670 290.205 ;
        RECT 3373.740 228.490 3374.000 228.810 ;
        RECT 3368.220 227.810 3368.480 228.130 ;
        RECT 3382.010 221.155 3382.290 221.525 ;
        RECT 2891.660 220.670 2891.920 220.990 ;
        RECT 2911.900 220.670 2912.160 220.990 ;
        RECT 2891.720 200.000 2891.860 220.670 ;
        RECT 3382.080 214.045 3382.220 221.155 ;
        RECT 3382.010 213.675 3382.290 214.045 ;
        RECT 2299.240 196.860 2319.285 198.000 ;
        RECT 2299.300 194.340 2319.285 196.860 ;
      LAYER met2 ;
        RECT 2319.565 197.395 2329.280 197.965 ;
      LAYER met2 ;
        RECT 2329.560 197.675 2339.560 198.000 ;
      LAYER met2 ;
        RECT 2339.840 197.395 2353.225 197.965 ;
        RECT 2319.565 196.235 2353.225 197.395 ;
      LAYER met2 ;
        RECT 2353.505 196.515 2373.500 198.000 ;
      LAYER met2 ;
        RECT 2319.565 194.060 2373.500 196.235 ;
        RECT 2299.300 3.570 2373.500 194.060 ;
      LAYER met2 ;
        RECT 2841.710 174.340 2865.610 200.000 ;
      LAYER met2 ;
        RECT 2865.890 197.665 2891.325 197.965 ;
      LAYER met2 ;
        RECT 2891.605 197.945 2915.505 200.000 ;
      LAYER met2 ;
        RECT 2865.890 174.060 2915.735 197.665 ;
        RECT 2841.710 4.925 2915.735 174.060 ;
      LAYER via2 ;
        RECT 1620.210 4982.560 1620.490 4982.840 ;
        RECT 200.650 4422.240 200.930 4422.520 ;
        RECT 200.650 4384.840 200.930 4385.120 ;
        RECT 210.770 4384.840 211.050 4385.120 ;
        RECT 223.190 4622.840 223.470 4623.120 ;
        RECT 224.110 4622.840 224.390 4623.120 ;
        RECT 386.490 4951.280 386.770 4951.560 ;
        RECT 414.090 4951.280 414.370 4951.560 ;
        RECT 510.690 4950.600 510.970 4950.880 ;
        RECT 531.390 4950.600 531.670 4950.880 ;
        RECT 966.090 4951.280 966.370 4951.560 ;
        RECT 1091.210 4951.280 1091.490 4951.560 ;
        RECT 1435.290 4952.640 1435.570 4952.920 ;
        RECT 1450.010 4952.640 1450.290 4952.920 ;
        RECT 2870.030 4985.280 2870.310 4985.560 ;
        RECT 1628.950 4952.640 1629.230 4952.920 ;
        RECT 1738.430 4952.640 1738.710 4952.920 ;
        RECT 1474.850 4951.280 1475.130 4951.560 ;
        RECT 1620.210 4951.280 1620.490 4951.560 ;
        RECT 223.190 4526.280 223.470 4526.560 ;
        RECT 224.110 4526.280 224.390 4526.560 ;
        RECT 223.650 4422.240 223.930 4422.520 ;
        RECT 220.890 4410.000 221.170 4410.280 ;
        RECT 224.110 4410.000 224.390 4410.280 ;
        RECT 223.650 4057.760 223.930 4058.040 ;
        RECT 223.190 4057.080 223.470 4057.360 ;
        RECT 3389.370 4405.920 3389.650 4406.200 ;
        RECT 3389.370 4380.760 3389.650 4381.040 ;
        RECT 223.190 3270.320 223.470 3270.600 ;
        RECT 224.110 3270.320 224.390 3270.600 ;
        RECT 211.230 2636.305 211.510 2636.585 ;
        RECT 223.190 2221.760 223.470 2222.040 ;
        RECT 224.110 2221.760 224.390 2222.040 ;
        RECT 3368.210 1958.600 3368.490 1958.880 ;
        RECT 223.650 1834.840 223.930 1835.120 ;
        RECT 224.110 1765.480 224.390 1765.760 ;
        RECT 3369.590 1932.080 3369.870 1932.360 ;
        RECT 223.650 773.360 223.930 773.640 ;
        RECT 223.190 772.680 223.470 772.960 ;
        RECT 224.110 385.760 224.390 386.040 ;
        RECT 224.110 289.880 224.390 290.160 ;
        RECT 676.290 202.160 676.570 202.440 ;
        RECT 1753.610 221.200 1753.890 221.480 ;
        RECT 1793.630 221.200 1793.910 221.480 ;
        RECT 741.150 200.800 741.430 201.080 ;
        RECT 1449.090 206.920 1449.370 207.200 ;
        RECT 1545.230 206.920 1545.510 207.200 ;
        RECT 1642.290 206.920 1642.570 207.200 ;
        RECT 1711.290 206.920 1711.570 207.200 ;
        RECT 1283.030 201.480 1283.310 201.760 ;
        RECT 717.690 198.080 717.970 198.360 ;
        RECT 2304.690 200.120 2304.970 200.400 ;
        RECT 2325.390 199.440 2325.670 199.720 ;
        RECT 2345.630 213.720 2345.910 214.000 ;
        RECT 2337.810 200.120 2338.090 200.400 ;
        RECT 2337.810 198.760 2338.090 199.040 ;
        RECT 2345.630 198.760 2345.910 199.040 ;
        RECT 3390.290 4363.760 3390.570 4364.040 ;
        RECT 3384.310 482.320 3384.590 482.600 ;
        RECT 3384.310 386.440 3384.590 386.720 ;
        RECT 3383.390 385.760 3383.670 386.040 ;
        RECT 3383.390 289.880 3383.670 290.160 ;
        RECT 3382.010 221.200 3382.290 221.480 ;
        RECT 3382.010 213.720 3382.290 214.000 ;
        RECT 2841.970 198.080 2842.250 198.360 ;
      LAYER met3 ;
        RECT 668.310 4986.690 747.570 5188.000 ;
        RECT 1213.310 4986.690 1292.570 5188.000 ;
        RECT 1758.310 4986.690 1837.570 5188.000 ;
        RECT 2303.310 4986.690 2382.570 5188.000 ;
        RECT 2848.240 5014.250 2922.290 5188.000 ;
      LAYER met3 ;
        RECT 2848.495 4988.000 2872.395 5013.850 ;
      LAYER met3 ;
        RECT 2872.795 5000.825 2897.990 5014.250 ;
        RECT 2872.795 5000.380 2873.495 5000.825 ;
        RECT 2885.295 5000.780 2897.990 5000.825 ;
      LAYER met3 ;
        RECT 2873.895 4988.000 2884.895 5000.425 ;
      LAYER met3 ;
        RECT 2885.295 5000.380 2885.490 5000.780 ;
        RECT 2897.290 5000.380 2897.990 5000.780 ;
      LAYER met3 ;
        RECT 2885.890 4988.000 2896.890 5000.380 ;
        RECT 2898.390 4988.000 2922.290 5013.850 ;
        RECT 2848.630 4985.570 2848.930 4988.000 ;
        RECT 2870.005 4985.570 2870.335 4985.585 ;
        RECT 2874.390 4985.570 2874.690 4988.000 ;
        RECT 2848.630 4985.270 2874.690 4985.570 ;
        RECT 2870.005 4985.255 2870.335 4985.270 ;
        RECT 1620.185 4982.850 1620.515 4982.865 ;
        RECT 2886.350 4982.850 2886.650 4988.000 ;
        RECT 1620.185 4982.550 2886.650 4982.850 ;
        RECT 1620.185 4982.535 1620.515 4982.550 ;
        RECT 1435.265 4952.930 1435.595 4952.945 ;
        RECT 1449.985 4952.930 1450.315 4952.945 ;
        RECT 1435.265 4952.630 1450.315 4952.930 ;
        RECT 1435.265 4952.615 1435.595 4952.630 ;
        RECT 1449.985 4952.615 1450.315 4952.630 ;
        RECT 1628.925 4952.930 1629.255 4952.945 ;
        RECT 1738.405 4952.930 1738.735 4952.945 ;
        RECT 1628.925 4952.630 1738.735 4952.930 ;
        RECT 1628.925 4952.615 1629.255 4952.630 ;
        RECT 1738.405 4952.615 1738.735 4952.630 ;
        RECT 386.465 4951.570 386.795 4951.585 ;
        RECT 414.065 4951.570 414.395 4951.585 ;
        RECT 386.465 4951.270 414.395 4951.570 ;
        RECT 386.465 4951.255 386.795 4951.270 ;
        RECT 414.065 4951.255 414.395 4951.270 ;
        RECT 966.065 4951.570 966.395 4951.585 ;
        RECT 1091.185 4951.570 1091.515 4951.585 ;
        RECT 966.065 4951.270 1091.515 4951.570 ;
        RECT 966.065 4951.255 966.395 4951.270 ;
        RECT 1091.185 4951.255 1091.515 4951.270 ;
        RECT 1474.825 4951.570 1475.155 4951.585 ;
        RECT 1620.185 4951.570 1620.515 4951.585 ;
        RECT 1474.825 4951.270 1620.515 4951.570 ;
        RECT 1474.825 4951.255 1475.155 4951.270 ;
        RECT 1620.185 4951.255 1620.515 4951.270 ;
        RECT 510.665 4950.890 510.995 4950.905 ;
        RECT 531.365 4950.890 531.695 4950.905 ;
        RECT 510.665 4950.590 531.695 4950.890 ;
        RECT 510.665 4950.575 510.995 4950.590 ;
        RECT 531.365 4950.575 531.695 4950.590 ;
        RECT 223.165 4623.130 223.495 4623.145 ;
        RECT 224.085 4623.130 224.415 4623.145 ;
        RECT 223.165 4622.830 224.415 4623.130 ;
        RECT 223.165 4622.815 223.495 4622.830 ;
        RECT 224.085 4622.815 224.415 4622.830 ;
        RECT 223.165 4526.570 223.495 4526.585 ;
        RECT 224.085 4526.570 224.415 4526.585 ;
        RECT 223.165 4526.270 224.415 4526.570 ;
        RECT 223.165 4526.255 223.495 4526.270 ;
        RECT 224.085 4526.255 224.415 4526.270 ;
      LAYER met3 ;
        RECT 0.000 4433.990 179.800 4458.290 ;
      LAYER met3 ;
        RECT 180.200 4434.390 200.000 4458.290 ;
      LAYER met3 ;
        RECT 0.000 4433.290 197.275 4433.990 ;
        RECT 0.000 4421.490 188.270 4433.290 ;
      LAYER met3 ;
        RECT 188.670 4422.530 200.000 4432.890 ;
        RECT 3390.000 4430.500 3396.900 4454.500 ;
      LAYER met3 ;
        RECT 3397.300 4430.100 3579.515 4454.510 ;
        RECT 3390.035 4429.400 3579.515 4430.100 ;
      LAYER met3 ;
        RECT 200.625 4422.530 200.955 4422.545 ;
        RECT 223.625 4422.530 223.955 4422.545 ;
        RECT 188.670 4422.230 223.955 4422.530 ;
        RECT 188.670 4421.890 200.000 4422.230 ;
        RECT 200.625 4422.215 200.955 4422.230 ;
        RECT 223.625 4422.215 223.955 4422.230 ;
      LAYER met3 ;
        RECT 0.000 4421.295 197.275 4421.490 ;
        RECT 0.000 4409.495 196.875 4421.295 ;
      LAYER met3 ;
        RECT 197.275 4410.290 200.000 4420.895 ;
        RECT 3390.000 4418.450 3410.220 4429.000 ;
        RECT 3388.670 4418.150 3410.220 4418.450 ;
        RECT 3388.670 4416.410 3388.970 4418.150 ;
        RECT 3390.000 4418.120 3410.220 4418.150 ;
      LAYER met3 ;
        RECT 3410.620 4417.720 3579.515 4429.400 ;
        RECT 3390.035 4417.020 3579.515 4417.720 ;
      LAYER met3 ;
        RECT 3390.000 4416.410 3412.900 4416.620 ;
        RECT 3388.670 4416.110 3412.900 4416.410 ;
        RECT 220.865 4410.290 221.195 4410.305 ;
        RECT 224.085 4410.290 224.415 4410.305 ;
        RECT 197.275 4409.990 224.415 4410.290 ;
        RECT 197.275 4409.895 200.000 4409.990 ;
        RECT 220.865 4409.975 221.195 4409.990 ;
        RECT 224.085 4409.975 224.415 4409.990 ;
      LAYER met3 ;
        RECT 0.000 4408.795 197.275 4409.495 ;
        RECT 0.000 4384.240 179.800 4408.795 ;
      LAYER met3 ;
        RECT 180.200 4385.130 200.000 4408.395 ;
        RECT 3389.345 4406.210 3389.675 4406.225 ;
        RECT 3390.000 4406.210 3412.900 4416.110 ;
        RECT 3389.345 4405.910 3412.900 4406.210 ;
        RECT 3389.345 4405.895 3389.675 4405.910 ;
        RECT 3390.000 4405.745 3412.900 4405.910 ;
      LAYER met3 ;
        RECT 3413.300 4405.345 3579.515 4417.020 ;
        RECT 3390.035 4404.645 3579.515 4405.345 ;
      LAYER met3 ;
        RECT 200.625 4385.130 200.955 4385.145 ;
        RECT 210.745 4385.130 211.075 4385.145 ;
        RECT 180.200 4384.830 211.075 4385.130 ;
        RECT 180.200 4384.495 200.000 4384.830 ;
        RECT 200.625 4384.815 200.955 4384.830 ;
        RECT 210.745 4384.815 211.075 4384.830 ;
        RECT 3389.345 4381.050 3389.675 4381.065 ;
        RECT 3390.000 4381.050 3396.900 4404.245 ;
        RECT 3389.345 4380.750 3396.900 4381.050 ;
        RECT 3389.345 4380.735 3389.675 4380.750 ;
        RECT 3390.000 4380.300 3396.900 4380.750 ;
      LAYER met3 ;
        RECT 3397.300 4380.300 3579.515 4404.645 ;
      LAYER met3 ;
        RECT 3387.710 4364.050 3388.090 4364.060 ;
        RECT 3390.265 4364.050 3390.595 4364.065 ;
        RECT 3387.710 4363.750 3390.595 4364.050 ;
        RECT 3387.710 4363.740 3388.090 4363.750 ;
        RECT 3390.265 4363.735 3390.595 4363.750 ;
        RECT 223.625 4058.050 223.955 4058.065 ;
        RECT 223.625 4057.735 224.170 4058.050 ;
        RECT 223.165 4057.370 223.495 4057.385 ;
        RECT 223.870 4057.370 224.170 4057.735 ;
        RECT 223.165 4057.070 224.170 4057.370 ;
        RECT 223.165 4057.055 223.495 4057.070 ;
      LAYER met3 ;
        RECT 0.000 3775.310 201.310 3854.570 ;
        RECT 3386.690 3771.430 3588.000 3850.690 ;
      LAYER met3 ;
        RECT 223.165 3270.610 223.495 3270.625 ;
        RECT 224.085 3270.610 224.415 3270.625 ;
        RECT 223.165 3270.310 224.415 3270.610 ;
        RECT 223.165 3270.295 223.495 3270.310 ;
        RECT 224.085 3270.295 224.415 3270.310 ;
      LAYER met3 ;
        RECT 0.000 3167.310 201.310 3246.570 ;
        RECT 3386.690 3163.430 3588.000 3242.690 ;
        RECT 0.000 2558.310 201.310 2637.570 ;
      LAYER met3 ;
        RECT 208.445 2636.595 208.775 2636.610 ;
        RECT 211.205 2636.595 211.535 2636.610 ;
        RECT 208.445 2636.295 211.535 2636.595 ;
        RECT 208.445 2636.280 208.775 2636.295 ;
        RECT 211.205 2636.280 211.535 2636.295 ;
      LAYER met3 ;
        RECT 3386.690 2554.430 3588.000 2633.690 ;
      LAYER met3 ;
        RECT 223.165 2222.050 223.495 2222.065 ;
        RECT 224.085 2222.050 224.415 2222.065 ;
        RECT 223.165 2221.750 224.415 2222.050 ;
        RECT 223.165 2221.735 223.495 2221.750 ;
        RECT 224.085 2221.735 224.415 2221.750 ;
      LAYER met3 ;
        RECT 0.000 1949.310 201.310 2028.570 ;
      LAYER met3 ;
        RECT 3368.185 1958.890 3368.515 1958.905 ;
        RECT 3369.310 1958.890 3369.690 1958.900 ;
        RECT 3368.185 1958.590 3369.690 1958.890 ;
        RECT 3368.185 1958.575 3368.515 1958.590 ;
        RECT 3369.310 1958.580 3369.690 1958.590 ;
      LAYER met3 ;
        RECT 3386.690 1945.430 3588.000 2024.690 ;
      LAYER met3 ;
        RECT 3369.565 1932.380 3369.895 1932.385 ;
        RECT 3369.310 1932.370 3369.895 1932.380 ;
        RECT 3369.310 1932.070 3370.120 1932.370 ;
        RECT 3369.310 1932.060 3369.895 1932.070 ;
        RECT 3369.565 1932.055 3369.895 1932.060 ;
        RECT 223.625 1835.140 223.955 1835.145 ;
        RECT 223.625 1835.130 224.210 1835.140 ;
        RECT 223.625 1834.830 224.410 1835.130 ;
        RECT 223.625 1834.820 224.210 1834.830 ;
        RECT 223.625 1834.815 223.955 1834.820 ;
        RECT 224.085 1765.780 224.415 1765.785 ;
        RECT 223.830 1765.770 224.415 1765.780 ;
        RECT 223.630 1765.470 224.415 1765.770 ;
        RECT 223.830 1765.460 224.415 1765.470 ;
        RECT 224.085 1765.455 224.415 1765.460 ;
      LAYER met3 ;
        RECT 0.000 1341.310 201.310 1420.570 ;
        RECT 3386.690 1337.430 3588.000 1416.690 ;
        RECT 0.000 732.310 201.310 811.570 ;
      LAYER met3 ;
        RECT 223.625 773.650 223.955 773.665 ;
        RECT 223.625 773.335 224.170 773.650 ;
        RECT 223.165 772.970 223.495 772.985 ;
        RECT 223.870 772.970 224.170 773.335 ;
        RECT 223.165 772.670 224.170 772.970 ;
        RECT 223.165 772.655 223.495 772.670 ;
      LAYER met3 ;
        RECT 3386.690 728.430 3588.000 807.690 ;
      LAYER met3 ;
        RECT 3381.270 510.490 3381.650 510.500 ;
        RECT 3384.950 510.490 3385.330 510.500 ;
        RECT 3381.270 510.190 3385.330 510.490 ;
        RECT 3381.270 510.180 3381.650 510.190 ;
        RECT 3384.950 510.180 3385.330 510.190 ;
        RECT 3384.285 482.610 3384.615 482.625 ;
        RECT 3384.950 482.610 3385.330 482.620 ;
        RECT 3384.285 482.310 3385.330 482.610 ;
        RECT 3384.285 482.295 3384.615 482.310 ;
        RECT 3384.950 482.300 3385.330 482.310 ;
        RECT 3384.285 386.740 3384.615 386.745 ;
        RECT 3384.030 386.730 3384.615 386.740 ;
        RECT 3383.830 386.430 3384.615 386.730 ;
        RECT 3384.030 386.420 3384.615 386.430 ;
        RECT 3384.285 386.415 3384.615 386.420 ;
        RECT 224.085 386.060 224.415 386.065 ;
        RECT 223.830 386.050 224.415 386.060 ;
        RECT 3383.365 386.050 3383.695 386.065 ;
        RECT 3384.030 386.050 3384.410 386.060 ;
        RECT 223.830 385.750 224.640 386.050 ;
        RECT 3383.365 385.750 3384.410 386.050 ;
        RECT 223.830 385.740 224.415 385.750 ;
        RECT 224.085 385.735 224.415 385.740 ;
        RECT 3383.365 385.735 3383.695 385.750 ;
        RECT 3384.030 385.740 3384.410 385.750 ;
        RECT 224.085 290.180 224.415 290.185 ;
        RECT 3383.365 290.180 3383.695 290.185 ;
        RECT 223.830 290.170 224.415 290.180 ;
        RECT 3383.110 290.170 3383.695 290.180 ;
        RECT 223.630 289.870 224.415 290.170 ;
        RECT 3382.910 289.870 3383.695 290.170 ;
        RECT 223.830 289.860 224.415 289.870 ;
        RECT 3383.110 289.860 3383.695 289.870 ;
        RECT 224.085 289.855 224.415 289.860 ;
        RECT 3383.365 289.855 3383.695 289.860 ;
        RECT 1753.585 221.490 1753.915 221.505 ;
        RECT 1793.605 221.490 1793.935 221.505 ;
        RECT 1753.585 221.190 1793.935 221.490 ;
        RECT 1753.585 221.175 1753.915 221.190 ;
        RECT 1793.605 221.175 1793.935 221.190 ;
        RECT 3381.985 221.490 3382.315 221.505 ;
        RECT 3383.110 221.490 3383.490 221.500 ;
        RECT 3381.985 221.190 3383.490 221.490 ;
        RECT 3381.985 221.175 3382.315 221.190 ;
        RECT 3383.110 221.180 3383.490 221.190 ;
        RECT 2345.605 214.010 2345.935 214.025 ;
        RECT 3381.985 214.010 3382.315 214.025 ;
        RECT 2345.605 213.710 3382.315 214.010 ;
        RECT 2345.605 213.695 2345.935 213.710 ;
        RECT 3381.985 213.695 3382.315 213.710 ;
        RECT 1449.065 207.210 1449.395 207.225 ;
        RECT 1545.205 207.210 1545.535 207.225 ;
        RECT 1449.065 206.910 1545.535 207.210 ;
        RECT 1449.065 206.895 1449.395 206.910 ;
        RECT 1545.205 206.895 1545.535 206.910 ;
        RECT 1642.265 207.210 1642.595 207.225 ;
        RECT 1711.265 207.210 1711.595 207.225 ;
        RECT 1642.265 206.910 1711.595 207.210 ;
        RECT 1642.265 206.895 1642.595 206.910 ;
        RECT 1711.265 206.895 1711.595 206.910 ;
        RECT 676.265 202.450 676.595 202.465 ;
        RECT 676.265 202.150 2842.490 202.450 ;
        RECT 676.265 202.135 676.595 202.150 ;
        RECT 1283.005 201.770 1283.335 201.785 ;
        RECT 1275.190 201.470 1283.335 201.770 ;
        RECT 741.125 201.090 741.455 201.105 ;
        RECT 717.910 200.790 741.455 201.090 ;
        RECT 717.910 200.000 718.210 200.790 ;
        RECT 741.125 200.775 741.455 200.790 ;
        RECT 1275.190 200.000 1275.490 201.470 ;
        RECT 1283.005 201.455 1283.335 201.470 ;
        RECT 667.710 163.240 691.610 200.000 ;
        RECT 693.110 187.620 704.110 200.000 ;
      LAYER met3 ;
        RECT 692.010 187.220 692.710 187.620 ;
        RECT 704.510 187.220 704.705 187.620 ;
      LAYER met3 ;
        RECT 705.105 187.575 716.105 200.000 ;
      LAYER met3 ;
        RECT 692.010 187.175 704.705 187.220 ;
        RECT 716.505 187.175 717.205 187.620 ;
        RECT 692.010 167.085 717.205 187.175 ;
      LAYER met3 ;
        RECT 717.605 167.485 741.505 200.000 ;
      LAYER met3 ;
        RECT 692.010 162.840 741.760 167.085 ;
        RECT 667.710 4.900 741.760 162.840 ;
        RECT 1209.300 151.080 1210.340 199.375 ;
        RECT 1209.300 133.400 1209.675 151.080 ;
      LAYER met3 ;
        RECT 1210.740 150.680 1211.810 200.000 ;
        RECT 1210.075 150.080 1211.810 150.680 ;
      LAYER met3 ;
        RECT 1212.210 188.690 1253.935 199.375 ;
        RECT 1255.465 193.730 1262.375 199.375 ;
        RECT 1255.465 192.265 1260.910 193.730 ;
      LAYER met3 ;
        RECT 1262.775 193.330 1263.925 200.000 ;
      LAYER met3 ;
        RECT 1255.465 191.985 1260.630 192.265 ;
      LAYER met3 ;
        RECT 1261.310 192.100 1263.925 193.330 ;
      LAYER met3 ;
        RECT 1255.465 190.555 1259.550 191.985 ;
      LAYER met3 ;
        RECT 1261.310 191.865 1262.775 192.100 ;
        RECT 1262.940 191.865 1263.925 192.100 ;
      LAYER met3 ;
        RECT 1264.325 196.465 1264.690 199.375 ;
      LAYER met3 ;
        RECT 1265.090 196.865 1266.755 200.000 ;
      LAYER met3 ;
        RECT 1267.155 196.465 1274.680 199.375 ;
      LAYER met3 ;
        RECT 1261.030 191.585 1261.310 191.865 ;
        RECT 1262.660 191.585 1262.940 191.865 ;
      LAYER met3 ;
        RECT 1255.765 190.255 1259.550 190.555 ;
        RECT 1212.210 184.830 1254.700 188.690 ;
        RECT 1256.230 187.335 1259.550 190.255 ;
      LAYER met3 ;
        RECT 1259.950 191.500 1261.030 191.585 ;
        RECT 1261.095 191.500 1262.660 191.585 ;
        RECT 1259.950 190.600 1262.660 191.500 ;
      LAYER met3 ;
        RECT 1264.325 191.465 1274.680 196.465 ;
        RECT 1263.340 191.185 1274.680 191.465 ;
      LAYER met3 ;
        RECT 1259.950 190.505 1261.030 190.600 ;
        RECT 1261.095 190.505 1262.660 190.600 ;
        RECT 1259.950 190.020 1262.660 190.505 ;
        RECT 1259.950 187.735 1261.095 190.020 ;
      LAYER met3 ;
        RECT 1263.060 189.620 1274.680 191.185 ;
        RECT 1261.495 187.335 1274.680 189.620 ;
        RECT 1256.230 184.830 1274.680 187.335 ;
        RECT 1212.210 183.015 1274.680 184.830 ;
      LAYER met3 ;
        RECT 1275.080 184.215 1275.600 200.000 ;
      LAYER met3 ;
        RECT 1276.000 184.615 1283.035 199.375 ;
        RECT 1276.210 184.405 1283.035 184.615 ;
      LAYER met3 ;
        RECT 1275.080 184.005 1275.810 184.215 ;
        RECT 1275.080 183.705 1275.670 184.005 ;
        RECT 1275.810 183.705 1276.260 184.005 ;
      LAYER met3 ;
        RECT 1276.660 183.955 1283.035 184.405 ;
      LAYER met3 ;
        RECT 1275.080 183.555 1276.260 183.705 ;
        RECT 1275.080 183.415 1275.670 183.555 ;
        RECT 1275.670 183.255 1276.130 183.415 ;
        RECT 1276.260 183.255 1276.710 183.555 ;
      LAYER met3 ;
        RECT 1277.110 183.505 1283.035 183.955 ;
      LAYER met3 ;
        RECT 1275.670 183.105 1276.710 183.255 ;
      LAYER met3 ;
        RECT 1212.210 182.555 1275.270 183.015 ;
      LAYER met3 ;
        RECT 1275.670 182.955 1277.225 183.105 ;
        RECT 1276.130 182.655 1276.705 182.955 ;
        RECT 1276.710 182.655 1277.225 182.955 ;
      LAYER met3 ;
        RECT 1212.210 181.980 1275.730 182.555 ;
      LAYER met3 ;
        RECT 1276.130 182.380 1277.225 182.655 ;
      LAYER met3 ;
        RECT 1212.210 169.105 1276.305 181.980 ;
        RECT 1212.210 168.520 1275.720 169.105 ;
      LAYER met3 ;
        RECT 1276.705 168.705 1277.225 182.380 ;
      LAYER met3 ;
        RECT 1212.210 167.805 1275.005 168.520 ;
      LAYER met3 ;
        RECT 1276.120 168.345 1277.225 168.705 ;
        RECT 1276.120 168.120 1276.705 168.345 ;
        RECT 1276.850 168.120 1277.225 168.345 ;
        RECT 1275.405 168.045 1276.120 168.120 ;
        RECT 1276.135 168.045 1276.850 168.120 ;
      LAYER met3 ;
        RECT 1212.210 167.220 1274.420 167.805 ;
      LAYER met3 ;
        RECT 1275.405 167.595 1276.850 168.045 ;
      LAYER met3 ;
        RECT 1277.625 167.720 1283.035 183.505 ;
      LAYER met3 ;
        RECT 1275.405 167.405 1276.120 167.595 ;
        RECT 1276.135 167.405 1276.850 167.595 ;
        RECT 1274.820 167.295 1275.405 167.405 ;
        RECT 1275.550 167.295 1276.135 167.405 ;
      LAYER met3 ;
        RECT 1212.210 167.005 1274.205 167.220 ;
        RECT 1212.210 165.475 1261.325 167.005 ;
      LAYER met3 ;
        RECT 1274.820 166.995 1276.135 167.295 ;
      LAYER met3 ;
        RECT 1277.250 167.005 1283.035 167.720 ;
      LAYER met3 ;
        RECT 1274.820 166.820 1275.405 166.995 ;
        RECT 1275.550 166.820 1276.135 166.995 ;
        RECT 1274.605 166.605 1274.820 166.820 ;
        RECT 1275.030 166.605 1275.550 166.820 ;
        RECT 1261.725 166.455 1275.550 166.605 ;
        RECT 1261.725 166.300 1274.885 166.305 ;
        RECT 1275.030 166.300 1275.550 166.455 ;
      LAYER met3 ;
        RECT 1276.535 166.420 1283.035 167.005 ;
      LAYER met3 ;
        RECT 1261.725 166.155 1275.030 166.300 ;
        RECT 1274.605 166.005 1275.030 166.155 ;
        RECT 1261.725 165.875 1275.030 166.005 ;
      LAYER met3 ;
        RECT 1275.950 165.900 1283.035 166.420 ;
        RECT 1275.430 165.475 1283.035 165.900 ;
      LAYER met3 ;
        RECT 1210.075 150.015 1210.740 150.080 ;
        RECT 1210.075 135.400 1211.810 150.015 ;
      LAYER met3 ;
        RECT 1212.210 135.800 1283.035 165.475 ;
      LAYER met3 ;
        RECT 1210.075 133.800 1213.410 135.400 ;
      LAYER met3 ;
        RECT 1213.810 134.200 1283.035 135.800 ;
        RECT 1209.300 131.800 1211.410 133.400 ;
      LAYER met3 ;
        RECT 1211.810 132.400 1214.810 133.800 ;
      LAYER met3 ;
        RECT 1215.210 132.800 1283.035 134.200 ;
      LAYER met3 ;
        RECT 1211.810 132.250 1215.745 132.400 ;
        RECT 1211.810 132.200 1213.410 132.250 ;
        RECT 1213.410 131.950 1214.695 132.200 ;
        RECT 1214.810 131.950 1215.745 132.250 ;
      LAYER met3 ;
        RECT 1209.300 130.515 1213.010 131.800 ;
      LAYER met3 ;
        RECT 1213.410 131.465 1215.745 131.950 ;
      LAYER met3 ;
        RECT 1216.145 131.865 1283.035 132.800 ;
      LAYER met3 ;
        RECT 1213.410 131.350 1215.710 131.465 ;
        RECT 1213.410 131.200 1214.695 131.350 ;
        RECT 1215.745 131.200 1216.610 131.465 ;
        RECT 1213.410 131.050 1216.610 131.200 ;
        RECT 1213.410 130.915 1214.695 131.050 ;
        RECT 1214.695 130.900 1215.645 130.915 ;
        RECT 1215.745 130.900 1216.610 131.050 ;
      LAYER met3 ;
        RECT 1217.010 131.000 1283.035 131.865 ;
      LAYER met3 ;
        RECT 1214.695 130.600 1216.610 130.900 ;
      LAYER met3 ;
        RECT 1209.300 129.565 1214.295 130.515 ;
      LAYER met3 ;
        RECT 1214.695 130.450 1217.960 130.600 ;
        RECT 1214.695 130.300 1215.645 130.450 ;
        RECT 1216.610 130.300 1217.960 130.450 ;
        RECT 1214.695 130.000 1217.960 130.300 ;
        RECT 1214.695 129.965 1215.645 130.000 ;
        RECT 1216.610 129.965 1217.960 130.000 ;
      LAYER met3 ;
        RECT 1209.300 128.600 1215.245 129.565 ;
      LAYER met3 ;
        RECT 1215.645 129.250 1217.960 129.965 ;
      LAYER met3 ;
        RECT 1218.360 129.650 1283.035 131.000 ;
      LAYER met3 ;
        RECT 1215.645 129.100 1219.140 129.250 ;
        RECT 1215.645 129.000 1216.610 129.100 ;
        RECT 1216.610 128.800 1217.820 129.000 ;
        RECT 1217.960 128.800 1219.140 129.100 ;
      LAYER met3 ;
        RECT 1209.300 127.390 1216.210 128.600 ;
      LAYER met3 ;
        RECT 1216.610 127.920 1219.140 128.800 ;
        RECT 1216.610 127.790 1217.820 127.920 ;
        RECT 1217.840 127.790 1219.140 127.920 ;
        RECT 1217.820 127.600 1219.140 127.790 ;
      LAYER met3 ;
        RECT 1209.300 127.200 1217.420 127.390 ;
        RECT 1209.300 104.955 1217.610 127.200 ;
      LAYER met3 ;
        RECT 1218.010 105.355 1219.140 127.600 ;
      LAYER met3 ;
        RECT 1219.540 104.955 1283.035 129.650 ;
        RECT 1209.300 0.000 1283.035 104.955 ;
        RECT 1752.430 0.000 1831.690 201.310 ;
      LAYER met3 ;
        RECT 2304.665 200.410 2304.995 200.425 ;
        RECT 2337.785 200.410 2338.115 200.425 ;
        RECT 2304.665 200.110 2338.115 200.410 ;
        RECT 2304.665 200.095 2304.995 200.110 ;
        RECT 2337.785 200.095 2338.115 200.110 ;
        RECT 2842.190 200.000 2842.490 202.150 ;
        RECT 2325.365 199.730 2325.695 199.745 ;
        RECT 2325.150 199.415 2325.695 199.730 ;
        RECT 2325.150 198.000 2325.450 199.415 ;
        RECT 2337.785 199.050 2338.115 199.065 ;
        RECT 2345.605 199.050 2345.935 199.065 ;
        RECT 2337.785 198.750 2350.290 199.050 ;
        RECT 2337.785 198.735 2338.115 198.750 ;
        RECT 2345.605 198.735 2345.935 198.750 ;
        RECT 2349.990 198.000 2350.290 198.750 ;
        RECT 2299.300 158.400 2323.245 198.000 ;
        RECT 2324.745 197.690 2335.620 198.000 ;
        RECT 2337.120 197.690 2348.000 198.000 ;
        RECT 2324.745 197.390 2348.000 197.690 ;
      LAYER met3 ;
        RECT 2323.645 174.700 2324.345 180.210 ;
      LAYER met3 ;
        RECT 2324.745 175.100 2335.620 197.390 ;
      LAYER met3 ;
        RECT 2336.020 177.380 2336.720 180.210 ;
      LAYER met3 ;
        RECT 2337.120 177.780 2348.000 197.390 ;
      LAYER met3 ;
        RECT 2348.400 177.380 2349.100 180.210 ;
        RECT 2336.020 174.700 2349.100 177.380 ;
        RECT 2323.645 158.000 2349.100 174.700 ;
      LAYER met3 ;
        RECT 2349.500 158.400 2373.500 198.000 ;
        RECT 2841.710 185.040 2865.610 200.000 ;
      LAYER met3 ;
        RECT 2866.010 188.270 2866.710 197.275 ;
      LAYER met3 ;
        RECT 2867.110 188.670 2878.110 200.000 ;
        RECT 2879.105 197.275 2890.105 200.000 ;
      LAYER met3 ;
        RECT 2878.510 196.875 2878.705 197.275 ;
        RECT 2890.505 196.875 2891.205 197.275 ;
        RECT 2878.510 188.270 2891.205 196.875 ;
        RECT 2866.010 184.640 2891.205 188.270 ;
      LAYER met3 ;
        RECT 2891.605 185.040 2915.505 200.000 ;
      LAYER met3 ;
        RECT 2299.300 8.485 2373.500 158.000 ;
        RECT 2841.345 0.000 2915.760 184.640 ;
      LAYER via3 ;
        RECT 3387.740 4363.740 3388.060 4364.060 ;
        RECT 3369.340 1958.580 3369.660 1958.900 ;
        RECT 3369.340 1932.060 3369.660 1932.380 ;
        RECT 223.860 1834.820 224.180 1835.140 ;
        RECT 223.860 1765.460 224.180 1765.780 ;
        RECT 3381.300 510.180 3381.620 510.500 ;
        RECT 3384.980 510.180 3385.300 510.500 ;
        RECT 3384.980 482.300 3385.300 482.620 ;
        RECT 3384.060 386.420 3384.380 386.740 ;
        RECT 223.860 385.740 224.180 386.060 ;
        RECT 3384.060 385.740 3384.380 386.060 ;
        RECT 223.860 289.860 224.180 290.180 ;
        RECT 3383.140 289.860 3383.460 290.180 ;
        RECT 3383.140 221.180 3383.460 221.500 ;
      LAYER met4 ;
        RECT 0.000 5163.385 202.330 5188.000 ;
      LAYER met4 ;
        RECT 202.730 5163.785 204.000 5188.000 ;
      LAYER met4 ;
        RECT 0.000 5083.400 202.745 5163.385 ;
        RECT 204.000 5162.035 668.000 5188.000 ;
      LAYER met4 ;
        RECT 668.000 5163.785 669.270 5188.000 ;
      LAYER met4 ;
        RECT 669.670 5163.385 746.330 5188.000 ;
      LAYER met4 ;
        RECT 746.730 5163.785 748.000 5188.000 ;
      LAYER met4 ;
        RECT 0.000 5057.635 201.745 5083.400 ;
        RECT 204.000 5083.000 668.000 5085.035 ;
        RECT 668.965 5083.400 746.970 5163.385 ;
        RECT 748.000 5162.035 1213.000 5188.000 ;
      LAYER met4 ;
        RECT 1213.000 5163.785 1214.270 5188.000 ;
      LAYER met4 ;
        RECT 1214.670 5163.385 1291.330 5188.000 ;
      LAYER met4 ;
        RECT 1291.730 5163.785 1293.000 5188.000 ;
        RECT 202.145 5058.035 205.000 5083.000 ;
      LAYER met4 ;
        RECT 205.000 5058.035 223.000 5083.000 ;
      LAYER met4 ;
        RECT 223.000 5058.035 225.000 5083.000 ;
      LAYER met4 ;
        RECT 225.000 5058.035 243.000 5083.000 ;
      LAYER met4 ;
        RECT 243.000 5058.035 245.000 5083.000 ;
      LAYER met4 ;
        RECT 245.000 5058.035 263.000 5083.000 ;
      LAYER met4 ;
        RECT 263.000 5058.035 265.000 5083.000 ;
      LAYER met4 ;
        RECT 265.000 5058.035 283.000 5083.000 ;
      LAYER met4 ;
        RECT 283.000 5058.035 285.000 5083.000 ;
      LAYER met4 ;
        RECT 285.000 5058.035 303.000 5083.000 ;
      LAYER met4 ;
        RECT 303.000 5058.035 305.000 5083.000 ;
      LAYER met4 ;
        RECT 305.000 5058.035 323.000 5083.000 ;
      LAYER met4 ;
        RECT 323.000 5058.035 325.000 5083.000 ;
      LAYER met4 ;
        RECT 325.000 5058.035 343.000 5083.000 ;
      LAYER met4 ;
        RECT 343.000 5058.035 345.000 5083.000 ;
      LAYER met4 ;
        RECT 345.000 5058.035 363.000 5083.000 ;
      LAYER met4 ;
        RECT 363.000 5058.035 365.000 5083.000 ;
      LAYER met4 ;
        RECT 365.000 5058.035 383.000 5083.000 ;
      LAYER met4 ;
        RECT 383.000 5058.035 385.000 5083.000 ;
      LAYER met4 ;
        RECT 385.000 5058.035 403.000 5083.000 ;
      LAYER met4 ;
        RECT 403.000 5058.035 405.000 5083.000 ;
      LAYER met4 ;
        RECT 405.000 5058.035 423.000 5083.000 ;
      LAYER met4 ;
        RECT 423.000 5058.035 425.000 5083.000 ;
      LAYER met4 ;
        RECT 425.000 5058.035 443.000 5083.000 ;
      LAYER met4 ;
        RECT 443.000 5058.035 445.000 5083.000 ;
      LAYER met4 ;
        RECT 445.000 5058.035 463.000 5083.000 ;
      LAYER met4 ;
        RECT 463.000 5058.035 465.000 5083.000 ;
      LAYER met4 ;
        RECT 465.000 5058.035 483.000 5083.000 ;
      LAYER met4 ;
        RECT 483.000 5058.035 485.000 5083.000 ;
      LAYER met4 ;
        RECT 485.000 5058.035 503.000 5083.000 ;
      LAYER met4 ;
        RECT 503.000 5058.035 505.000 5083.000 ;
      LAYER met4 ;
        RECT 505.000 5058.035 523.000 5083.000 ;
      LAYER met4 ;
        RECT 523.000 5058.035 525.000 5083.000 ;
      LAYER met4 ;
        RECT 525.000 5058.035 543.000 5083.000 ;
      LAYER met4 ;
        RECT 543.000 5058.035 545.000 5083.000 ;
      LAYER met4 ;
        RECT 545.000 5058.035 563.000 5083.000 ;
      LAYER met4 ;
        RECT 563.000 5058.035 565.000 5083.000 ;
      LAYER met4 ;
        RECT 565.000 5058.035 583.000 5083.000 ;
      LAYER met4 ;
        RECT 583.000 5058.035 585.000 5083.000 ;
      LAYER met4 ;
        RECT 585.000 5058.035 603.000 5083.000 ;
      LAYER met4 ;
        RECT 603.000 5058.035 605.000 5083.000 ;
      LAYER met4 ;
        RECT 605.000 5058.035 623.000 5083.000 ;
      LAYER met4 ;
        RECT 623.000 5058.035 625.000 5083.000 ;
      LAYER met4 ;
        RECT 625.000 5058.035 643.000 5083.000 ;
      LAYER met4 ;
        RECT 643.000 5058.035 645.000 5083.000 ;
      LAYER met4 ;
        RECT 645.000 5058.035 663.000 5083.000 ;
      LAYER met4 ;
        RECT 663.000 5058.035 669.270 5083.000 ;
      LAYER met4 ;
        RECT 0.000 5056.935 202.745 5057.635 ;
        RECT 204.000 5056.935 668.000 5058.035 ;
        RECT 669.670 5057.635 746.330 5083.400 ;
        RECT 748.000 5083.000 1213.000 5085.035 ;
        RECT 1213.965 5083.400 1291.970 5163.385 ;
        RECT 1293.000 5162.035 1758.000 5188.000 ;
      LAYER met4 ;
        RECT 1758.000 5163.785 1759.270 5188.000 ;
      LAYER met4 ;
        RECT 1759.670 5163.385 1836.330 5188.000 ;
      LAYER met4 ;
        RECT 1836.730 5163.785 1838.000 5188.000 ;
        RECT 746.730 5058.035 749.000 5083.000 ;
      LAYER met4 ;
        RECT 749.000 5058.035 767.000 5083.000 ;
      LAYER met4 ;
        RECT 767.000 5058.035 769.000 5083.000 ;
      LAYER met4 ;
        RECT 769.000 5058.035 787.000 5083.000 ;
      LAYER met4 ;
        RECT 787.000 5058.035 789.000 5083.000 ;
      LAYER met4 ;
        RECT 789.000 5058.035 807.000 5083.000 ;
      LAYER met4 ;
        RECT 807.000 5058.035 809.000 5083.000 ;
      LAYER met4 ;
        RECT 809.000 5058.035 827.000 5083.000 ;
      LAYER met4 ;
        RECT 827.000 5058.035 829.000 5083.000 ;
      LAYER met4 ;
        RECT 829.000 5058.035 847.000 5083.000 ;
      LAYER met4 ;
        RECT 847.000 5058.035 849.000 5083.000 ;
      LAYER met4 ;
        RECT 849.000 5058.035 867.000 5083.000 ;
      LAYER met4 ;
        RECT 867.000 5058.035 869.000 5083.000 ;
      LAYER met4 ;
        RECT 869.000 5058.035 887.000 5083.000 ;
      LAYER met4 ;
        RECT 887.000 5058.035 889.000 5083.000 ;
      LAYER met4 ;
        RECT 889.000 5058.035 907.000 5083.000 ;
      LAYER met4 ;
        RECT 907.000 5058.035 909.000 5083.000 ;
      LAYER met4 ;
        RECT 909.000 5058.035 927.000 5083.000 ;
      LAYER met4 ;
        RECT 927.000 5058.035 929.000 5083.000 ;
      LAYER met4 ;
        RECT 929.000 5058.035 947.000 5083.000 ;
      LAYER met4 ;
        RECT 947.000 5058.035 949.000 5083.000 ;
      LAYER met4 ;
        RECT 949.000 5058.035 967.000 5083.000 ;
      LAYER met4 ;
        RECT 967.000 5058.035 969.000 5083.000 ;
      LAYER met4 ;
        RECT 969.000 5058.035 987.000 5083.000 ;
      LAYER met4 ;
        RECT 987.000 5058.035 989.000 5083.000 ;
      LAYER met4 ;
        RECT 989.000 5058.035 1007.000 5083.000 ;
      LAYER met4 ;
        RECT 1007.000 5058.035 1009.000 5083.000 ;
      LAYER met4 ;
        RECT 1009.000 5058.035 1027.000 5083.000 ;
      LAYER met4 ;
        RECT 1027.000 5058.035 1029.000 5083.000 ;
      LAYER met4 ;
        RECT 1029.000 5058.035 1047.000 5083.000 ;
      LAYER met4 ;
        RECT 1047.000 5058.035 1049.000 5083.000 ;
      LAYER met4 ;
        RECT 1049.000 5058.035 1067.000 5083.000 ;
      LAYER met4 ;
        RECT 1067.000 5058.035 1069.000 5083.000 ;
      LAYER met4 ;
        RECT 1069.000 5058.035 1087.000 5083.000 ;
      LAYER met4 ;
        RECT 1087.000 5058.035 1089.000 5083.000 ;
      LAYER met4 ;
        RECT 1089.000 5058.035 1107.000 5083.000 ;
      LAYER met4 ;
        RECT 1107.000 5058.035 1109.000 5083.000 ;
      LAYER met4 ;
        RECT 1109.000 5058.035 1127.000 5083.000 ;
      LAYER met4 ;
        RECT 1127.000 5058.035 1129.000 5083.000 ;
      LAYER met4 ;
        RECT 1129.000 5058.035 1147.000 5083.000 ;
      LAYER met4 ;
        RECT 1147.000 5058.035 1149.000 5083.000 ;
      LAYER met4 ;
        RECT 1149.000 5058.035 1167.000 5083.000 ;
      LAYER met4 ;
        RECT 1167.000 5058.035 1169.000 5083.000 ;
      LAYER met4 ;
        RECT 1169.000 5058.035 1187.000 5083.000 ;
      LAYER met4 ;
        RECT 1187.000 5058.035 1189.000 5083.000 ;
      LAYER met4 ;
        RECT 1189.000 5058.035 1207.000 5083.000 ;
      LAYER met4 ;
        RECT 1207.000 5058.035 1209.000 5083.000 ;
      LAYER met4 ;
        RECT 1209.000 5058.035 1212.000 5083.000 ;
      LAYER met4 ;
        RECT 1212.000 5058.035 1214.270 5083.000 ;
      LAYER met4 ;
        RECT 668.965 5056.935 746.970 5057.635 ;
        RECT 748.000 5056.935 1213.000 5058.035 ;
        RECT 1214.670 5057.635 1291.330 5083.400 ;
        RECT 1293.000 5083.000 1758.000 5085.035 ;
        RECT 1758.965 5083.400 1836.970 5163.385 ;
        RECT 1838.000 5162.035 2303.000 5188.000 ;
      LAYER met4 ;
        RECT 2303.000 5163.785 2304.270 5188.000 ;
      LAYER met4 ;
        RECT 2304.670 5163.385 2381.330 5188.000 ;
      LAYER met4 ;
        RECT 2381.730 5163.785 2383.000 5188.000 ;
        RECT 1291.730 5058.035 1294.000 5083.000 ;
      LAYER met4 ;
        RECT 1294.000 5058.035 1312.000 5083.000 ;
      LAYER met4 ;
        RECT 1312.000 5058.035 1314.000 5083.000 ;
      LAYER met4 ;
        RECT 1314.000 5058.035 1332.000 5083.000 ;
      LAYER met4 ;
        RECT 1332.000 5058.035 1334.000 5083.000 ;
      LAYER met4 ;
        RECT 1334.000 5058.035 1352.000 5083.000 ;
      LAYER met4 ;
        RECT 1352.000 5058.035 1354.000 5083.000 ;
      LAYER met4 ;
        RECT 1354.000 5058.035 1372.000 5083.000 ;
      LAYER met4 ;
        RECT 1372.000 5058.035 1374.000 5083.000 ;
      LAYER met4 ;
        RECT 1374.000 5058.035 1392.000 5083.000 ;
      LAYER met4 ;
        RECT 1392.000 5058.035 1394.000 5083.000 ;
      LAYER met4 ;
        RECT 1394.000 5058.035 1412.000 5083.000 ;
      LAYER met4 ;
        RECT 1412.000 5058.035 1414.000 5083.000 ;
      LAYER met4 ;
        RECT 1414.000 5058.035 1432.000 5083.000 ;
      LAYER met4 ;
        RECT 1432.000 5058.035 1434.000 5083.000 ;
      LAYER met4 ;
        RECT 1434.000 5058.035 1452.000 5083.000 ;
      LAYER met4 ;
        RECT 1452.000 5058.035 1454.000 5083.000 ;
      LAYER met4 ;
        RECT 1454.000 5058.035 1472.000 5083.000 ;
      LAYER met4 ;
        RECT 1472.000 5058.035 1474.000 5083.000 ;
      LAYER met4 ;
        RECT 1474.000 5058.035 1492.000 5083.000 ;
      LAYER met4 ;
        RECT 1492.000 5058.035 1494.000 5083.000 ;
      LAYER met4 ;
        RECT 1494.000 5058.035 1512.000 5083.000 ;
      LAYER met4 ;
        RECT 1512.000 5058.035 1514.000 5083.000 ;
      LAYER met4 ;
        RECT 1514.000 5058.035 1532.000 5083.000 ;
      LAYER met4 ;
        RECT 1532.000 5058.035 1534.000 5083.000 ;
      LAYER met4 ;
        RECT 1534.000 5058.035 1552.000 5083.000 ;
      LAYER met4 ;
        RECT 1552.000 5058.035 1554.000 5083.000 ;
      LAYER met4 ;
        RECT 1554.000 5058.035 1572.000 5083.000 ;
      LAYER met4 ;
        RECT 1572.000 5058.035 1574.000 5083.000 ;
      LAYER met4 ;
        RECT 1574.000 5058.035 1592.000 5083.000 ;
      LAYER met4 ;
        RECT 1592.000 5058.035 1594.000 5083.000 ;
      LAYER met4 ;
        RECT 1594.000 5058.035 1612.000 5083.000 ;
      LAYER met4 ;
        RECT 1612.000 5058.035 1614.000 5083.000 ;
      LAYER met4 ;
        RECT 1614.000 5058.035 1632.000 5083.000 ;
      LAYER met4 ;
        RECT 1632.000 5058.035 1634.000 5083.000 ;
      LAYER met4 ;
        RECT 1634.000 5058.035 1652.000 5083.000 ;
      LAYER met4 ;
        RECT 1652.000 5058.035 1654.000 5083.000 ;
      LAYER met4 ;
        RECT 1654.000 5058.035 1672.000 5083.000 ;
      LAYER met4 ;
        RECT 1672.000 5058.035 1674.000 5083.000 ;
      LAYER met4 ;
        RECT 1674.000 5058.035 1692.000 5083.000 ;
      LAYER met4 ;
        RECT 1692.000 5058.035 1694.000 5083.000 ;
      LAYER met4 ;
        RECT 1694.000 5058.035 1712.000 5083.000 ;
      LAYER met4 ;
        RECT 1712.000 5058.035 1714.000 5083.000 ;
      LAYER met4 ;
        RECT 1714.000 5058.035 1732.000 5083.000 ;
      LAYER met4 ;
        RECT 1732.000 5058.035 1734.000 5083.000 ;
      LAYER met4 ;
        RECT 1734.000 5058.035 1752.000 5083.000 ;
      LAYER met4 ;
        RECT 1752.000 5058.035 1754.000 5083.000 ;
      LAYER met4 ;
        RECT 1754.000 5058.035 1757.000 5083.000 ;
      LAYER met4 ;
        RECT 1757.000 5058.035 1759.270 5083.000 ;
      LAYER met4 ;
        RECT 1213.965 5056.935 1291.970 5057.635 ;
        RECT 1293.000 5056.935 1758.000 5058.035 ;
        RECT 1759.670 5057.635 1836.330 5083.400 ;
        RECT 1838.000 5083.000 2303.000 5085.035 ;
        RECT 2303.965 5083.400 2381.970 5163.385 ;
        RECT 2383.000 5162.035 2848.000 5188.000 ;
      LAYER met4 ;
        RECT 2848.000 5163.785 2849.270 5188.000 ;
      LAYER met4 ;
        RECT 2849.670 5163.385 2921.330 5188.000 ;
      LAYER met4 ;
        RECT 2921.730 5163.785 2923.000 5188.000 ;
      LAYER met4 ;
        RECT 2923.000 5163.385 3388.000 5188.000 ;
      LAYER met4 ;
        RECT 3388.000 5163.785 3389.435 5188.000 ;
      LAYER met4 ;
        RECT 3389.835 5163.385 3588.000 5188.000 ;
      LAYER met4 ;
        RECT 1836.730 5058.035 1839.000 5083.000 ;
      LAYER met4 ;
        RECT 1839.000 5058.035 1857.000 5083.000 ;
      LAYER met4 ;
        RECT 1857.000 5058.035 1859.000 5083.000 ;
      LAYER met4 ;
        RECT 1859.000 5058.035 1877.000 5083.000 ;
      LAYER met4 ;
        RECT 1877.000 5058.035 1879.000 5083.000 ;
      LAYER met4 ;
        RECT 1879.000 5058.035 1897.000 5083.000 ;
      LAYER met4 ;
        RECT 1897.000 5058.035 1899.000 5083.000 ;
      LAYER met4 ;
        RECT 1899.000 5058.035 1917.000 5083.000 ;
      LAYER met4 ;
        RECT 1917.000 5058.035 1919.000 5083.000 ;
      LAYER met4 ;
        RECT 1919.000 5058.035 1937.000 5083.000 ;
      LAYER met4 ;
        RECT 1937.000 5058.035 1939.000 5083.000 ;
      LAYER met4 ;
        RECT 1939.000 5058.035 1957.000 5083.000 ;
      LAYER met4 ;
        RECT 1957.000 5058.035 1959.000 5083.000 ;
      LAYER met4 ;
        RECT 1959.000 5058.035 1977.000 5083.000 ;
      LAYER met4 ;
        RECT 1977.000 5058.035 1979.000 5083.000 ;
      LAYER met4 ;
        RECT 1979.000 5058.035 1997.000 5083.000 ;
      LAYER met4 ;
        RECT 1997.000 5058.035 1999.000 5083.000 ;
      LAYER met4 ;
        RECT 1999.000 5058.035 2017.000 5083.000 ;
      LAYER met4 ;
        RECT 2017.000 5058.035 2019.000 5083.000 ;
      LAYER met4 ;
        RECT 2019.000 5058.035 2037.000 5083.000 ;
      LAYER met4 ;
        RECT 2037.000 5058.035 2039.000 5083.000 ;
      LAYER met4 ;
        RECT 2039.000 5058.035 2057.000 5083.000 ;
      LAYER met4 ;
        RECT 2057.000 5058.035 2059.000 5083.000 ;
      LAYER met4 ;
        RECT 2059.000 5058.035 2077.000 5083.000 ;
      LAYER met4 ;
        RECT 2077.000 5058.035 2079.000 5083.000 ;
      LAYER met4 ;
        RECT 2079.000 5058.035 2097.000 5083.000 ;
      LAYER met4 ;
        RECT 2097.000 5058.035 2099.000 5083.000 ;
      LAYER met4 ;
        RECT 2099.000 5058.035 2117.000 5083.000 ;
      LAYER met4 ;
        RECT 2117.000 5058.035 2119.000 5083.000 ;
      LAYER met4 ;
        RECT 2119.000 5058.035 2137.000 5083.000 ;
      LAYER met4 ;
        RECT 2137.000 5058.035 2139.000 5083.000 ;
      LAYER met4 ;
        RECT 2139.000 5058.035 2157.000 5083.000 ;
      LAYER met4 ;
        RECT 2157.000 5058.035 2159.000 5083.000 ;
      LAYER met4 ;
        RECT 2159.000 5058.035 2177.000 5083.000 ;
      LAYER met4 ;
        RECT 2177.000 5058.035 2179.000 5083.000 ;
      LAYER met4 ;
        RECT 2179.000 5058.035 2197.000 5083.000 ;
      LAYER met4 ;
        RECT 2197.000 5058.035 2199.000 5083.000 ;
      LAYER met4 ;
        RECT 2199.000 5058.035 2217.000 5083.000 ;
      LAYER met4 ;
        RECT 2217.000 5058.035 2219.000 5083.000 ;
      LAYER met4 ;
        RECT 2219.000 5058.035 2237.000 5083.000 ;
      LAYER met4 ;
        RECT 2237.000 5058.035 2239.000 5083.000 ;
      LAYER met4 ;
        RECT 2239.000 5058.035 2257.000 5083.000 ;
      LAYER met4 ;
        RECT 2257.000 5058.035 2259.000 5083.000 ;
      LAYER met4 ;
        RECT 2259.000 5058.035 2277.000 5083.000 ;
      LAYER met4 ;
        RECT 2277.000 5058.035 2279.000 5083.000 ;
      LAYER met4 ;
        RECT 2279.000 5058.035 2297.000 5083.000 ;
      LAYER met4 ;
        RECT 2297.000 5058.035 2299.000 5083.000 ;
      LAYER met4 ;
        RECT 2299.000 5058.035 2302.000 5083.000 ;
      LAYER met4 ;
        RECT 2302.000 5058.035 2304.270 5083.000 ;
      LAYER met4 ;
        RECT 1758.965 5056.935 1836.970 5057.635 ;
        RECT 1838.000 5056.935 2303.000 5058.035 ;
        RECT 2304.670 5057.635 2381.330 5083.400 ;
        RECT 2383.000 5083.000 2848.000 5085.035 ;
        RECT 2848.965 5083.400 2922.035 5163.385 ;
        RECT 2923.000 5162.035 3588.000 5163.385 ;
        RECT 3388.000 5085.035 3588.000 5162.035 ;
        RECT 2923.000 5083.400 3588.000 5085.035 ;
      LAYER met4 ;
        RECT 2381.730 5058.035 2384.000 5083.000 ;
      LAYER met4 ;
        RECT 2384.000 5058.035 2402.000 5083.000 ;
      LAYER met4 ;
        RECT 2402.000 5058.035 2404.000 5083.000 ;
      LAYER met4 ;
        RECT 2404.000 5058.035 2422.000 5083.000 ;
      LAYER met4 ;
        RECT 2422.000 5058.035 2424.000 5083.000 ;
      LAYER met4 ;
        RECT 2424.000 5058.035 2442.000 5083.000 ;
      LAYER met4 ;
        RECT 2442.000 5058.035 2444.000 5083.000 ;
      LAYER met4 ;
        RECT 2444.000 5058.035 2462.000 5083.000 ;
      LAYER met4 ;
        RECT 2462.000 5058.035 2464.000 5083.000 ;
      LAYER met4 ;
        RECT 2464.000 5058.035 2482.000 5083.000 ;
      LAYER met4 ;
        RECT 2482.000 5058.035 2484.000 5083.000 ;
      LAYER met4 ;
        RECT 2484.000 5058.035 2502.000 5083.000 ;
      LAYER met4 ;
        RECT 2502.000 5058.035 2504.000 5083.000 ;
      LAYER met4 ;
        RECT 2504.000 5058.035 2522.000 5083.000 ;
      LAYER met4 ;
        RECT 2522.000 5058.035 2524.000 5083.000 ;
      LAYER met4 ;
        RECT 2524.000 5058.035 2542.000 5083.000 ;
      LAYER met4 ;
        RECT 2542.000 5058.035 2544.000 5083.000 ;
      LAYER met4 ;
        RECT 2544.000 5058.035 2562.000 5083.000 ;
      LAYER met4 ;
        RECT 2562.000 5058.035 2564.000 5083.000 ;
      LAYER met4 ;
        RECT 2564.000 5058.035 2582.000 5083.000 ;
      LAYER met4 ;
        RECT 2582.000 5058.035 2584.000 5083.000 ;
      LAYER met4 ;
        RECT 2584.000 5058.035 2602.000 5083.000 ;
      LAYER met4 ;
        RECT 2602.000 5058.035 2604.000 5083.000 ;
      LAYER met4 ;
        RECT 2604.000 5058.035 2622.000 5083.000 ;
      LAYER met4 ;
        RECT 2622.000 5058.035 2624.000 5083.000 ;
      LAYER met4 ;
        RECT 2624.000 5058.035 2642.000 5083.000 ;
      LAYER met4 ;
        RECT 2642.000 5058.035 2644.000 5083.000 ;
      LAYER met4 ;
        RECT 2644.000 5058.035 2662.000 5083.000 ;
      LAYER met4 ;
        RECT 2662.000 5058.035 2664.000 5083.000 ;
      LAYER met4 ;
        RECT 2664.000 5058.035 2682.000 5083.000 ;
      LAYER met4 ;
        RECT 2682.000 5058.035 2684.000 5083.000 ;
      LAYER met4 ;
        RECT 2684.000 5058.035 2702.000 5083.000 ;
      LAYER met4 ;
        RECT 2702.000 5058.035 2704.000 5083.000 ;
      LAYER met4 ;
        RECT 2704.000 5058.035 2722.000 5083.000 ;
      LAYER met4 ;
        RECT 2722.000 5058.035 2724.000 5083.000 ;
      LAYER met4 ;
        RECT 2724.000 5058.035 2742.000 5083.000 ;
      LAYER met4 ;
        RECT 2742.000 5058.035 2744.000 5083.000 ;
      LAYER met4 ;
        RECT 2744.000 5058.035 2762.000 5083.000 ;
      LAYER met4 ;
        RECT 2762.000 5058.035 2764.000 5083.000 ;
      LAYER met4 ;
        RECT 2764.000 5058.035 2782.000 5083.000 ;
      LAYER met4 ;
        RECT 2782.000 5058.035 2784.000 5083.000 ;
      LAYER met4 ;
        RECT 2784.000 5058.035 2802.000 5083.000 ;
      LAYER met4 ;
        RECT 2802.000 5058.035 2804.000 5083.000 ;
      LAYER met4 ;
        RECT 2804.000 5058.035 2822.000 5083.000 ;
      LAYER met4 ;
        RECT 2822.000 5058.035 2824.000 5083.000 ;
      LAYER met4 ;
        RECT 2824.000 5058.035 2842.000 5083.000 ;
      LAYER met4 ;
        RECT 2842.000 5058.035 2844.000 5083.000 ;
      LAYER met4 ;
        RECT 2844.000 5058.035 2847.000 5083.000 ;
      LAYER met4 ;
        RECT 2847.000 5058.035 2849.270 5083.000 ;
      LAYER met4 ;
        RECT 2303.965 5056.935 2381.970 5057.635 ;
        RECT 2383.000 5056.935 2848.000 5058.035 ;
        RECT 2849.670 5057.635 2921.330 5083.400 ;
        RECT 2923.000 5083.000 3388.000 5083.400 ;
      LAYER met4 ;
        RECT 2921.730 5058.035 2924.000 5083.000 ;
      LAYER met4 ;
        RECT 2924.000 5058.035 2942.000 5083.000 ;
      LAYER met4 ;
        RECT 2942.000 5058.035 2944.000 5083.000 ;
      LAYER met4 ;
        RECT 2944.000 5058.035 2962.000 5083.000 ;
      LAYER met4 ;
        RECT 2962.000 5058.035 2964.000 5083.000 ;
      LAYER met4 ;
        RECT 2964.000 5058.035 2982.000 5083.000 ;
      LAYER met4 ;
        RECT 2982.000 5058.035 2984.000 5083.000 ;
      LAYER met4 ;
        RECT 2984.000 5058.035 3002.000 5083.000 ;
      LAYER met4 ;
        RECT 3002.000 5058.035 3004.000 5083.000 ;
      LAYER met4 ;
        RECT 3004.000 5058.035 3022.000 5083.000 ;
      LAYER met4 ;
        RECT 3022.000 5058.035 3024.000 5083.000 ;
      LAYER met4 ;
        RECT 3024.000 5058.035 3042.000 5083.000 ;
      LAYER met4 ;
        RECT 3042.000 5058.035 3044.000 5083.000 ;
      LAYER met4 ;
        RECT 3044.000 5058.035 3062.000 5083.000 ;
      LAYER met4 ;
        RECT 3062.000 5058.035 3064.000 5083.000 ;
      LAYER met4 ;
        RECT 3064.000 5058.035 3082.000 5083.000 ;
      LAYER met4 ;
        RECT 3082.000 5058.035 3084.000 5083.000 ;
      LAYER met4 ;
        RECT 3084.000 5058.035 3102.000 5083.000 ;
      LAYER met4 ;
        RECT 3102.000 5058.035 3104.000 5083.000 ;
      LAYER met4 ;
        RECT 3104.000 5058.035 3122.000 5083.000 ;
      LAYER met4 ;
        RECT 3122.000 5058.035 3124.000 5083.000 ;
      LAYER met4 ;
        RECT 3124.000 5058.035 3142.000 5083.000 ;
      LAYER met4 ;
        RECT 3142.000 5058.035 3144.000 5083.000 ;
      LAYER met4 ;
        RECT 3144.000 5058.035 3162.000 5083.000 ;
      LAYER met4 ;
        RECT 3162.000 5058.035 3164.000 5083.000 ;
      LAYER met4 ;
        RECT 3164.000 5058.035 3182.000 5083.000 ;
      LAYER met4 ;
        RECT 3182.000 5058.035 3184.000 5083.000 ;
      LAYER met4 ;
        RECT 3184.000 5058.035 3202.000 5083.000 ;
      LAYER met4 ;
        RECT 3202.000 5058.035 3204.000 5083.000 ;
      LAYER met4 ;
        RECT 3204.000 5058.035 3222.000 5083.000 ;
      LAYER met4 ;
        RECT 3222.000 5058.035 3224.000 5083.000 ;
      LAYER met4 ;
        RECT 3224.000 5058.035 3242.000 5083.000 ;
      LAYER met4 ;
        RECT 3242.000 5058.035 3244.000 5083.000 ;
      LAYER met4 ;
        RECT 3244.000 5058.035 3262.000 5083.000 ;
      LAYER met4 ;
        RECT 3262.000 5058.035 3264.000 5083.000 ;
      LAYER met4 ;
        RECT 3264.000 5058.035 3282.000 5083.000 ;
      LAYER met4 ;
        RECT 3282.000 5058.035 3284.000 5083.000 ;
      LAYER met4 ;
        RECT 3284.000 5058.035 3302.000 5083.000 ;
      LAYER met4 ;
        RECT 3302.000 5058.035 3304.000 5083.000 ;
      LAYER met4 ;
        RECT 3304.000 5058.035 3322.000 5083.000 ;
      LAYER met4 ;
        RECT 3322.000 5058.035 3324.000 5083.000 ;
      LAYER met4 ;
        RECT 3324.000 5058.035 3342.000 5083.000 ;
      LAYER met4 ;
        RECT 3342.000 5058.035 3344.000 5083.000 ;
      LAYER met4 ;
        RECT 3344.000 5058.035 3362.000 5083.000 ;
      LAYER met4 ;
        RECT 3362.000 5058.035 3364.000 5083.000 ;
      LAYER met4 ;
        RECT 3364.000 5058.035 3382.000 5083.000 ;
      LAYER met4 ;
        RECT 3382.000 5058.035 3384.000 5083.000 ;
      LAYER met4 ;
        RECT 3384.000 5058.035 3387.000 5083.000 ;
      LAYER met4 ;
        RECT 3387.000 5058.035 3390.645 5083.000 ;
      LAYER met4 ;
        RECT 2923.000 5057.635 3388.000 5058.035 ;
        RECT 3391.045 5057.635 3588.000 5083.400 ;
        RECT 2848.965 5056.935 2922.035 5057.635 ;
        RECT 2923.000 5056.935 3588.000 5057.635 ;
        RECT 0.000 5051.685 202.330 5056.935 ;
      LAYER met4 ;
        RECT 202.730 5052.085 669.270 5056.535 ;
      LAYER met4 ;
        RECT 669.670 5051.685 746.330 5056.935 ;
      LAYER met4 ;
        RECT 746.730 5052.085 1214.270 5056.535 ;
      LAYER met4 ;
        RECT 1214.670 5051.685 1291.330 5056.935 ;
      LAYER met4 ;
        RECT 1291.730 5052.085 1759.270 5056.535 ;
      LAYER met4 ;
        RECT 1759.670 5051.685 1836.330 5056.935 ;
      LAYER met4 ;
        RECT 1836.730 5052.085 2304.270 5056.535 ;
      LAYER met4 ;
        RECT 2304.670 5051.685 2381.330 5056.935 ;
      LAYER met4 ;
        RECT 2381.730 5052.085 2849.270 5056.535 ;
      LAYER met4 ;
        RECT 2849.670 5051.685 2921.330 5056.935 ;
      LAYER met4 ;
        RECT 2921.730 5052.085 3389.480 5056.535 ;
      LAYER met4 ;
        RECT 3389.880 5051.685 3588.000 5056.935 ;
        RECT 0.000 5051.085 202.745 5051.685 ;
        RECT 204.000 5051.085 664.000 5051.685 ;
        RECT 668.965 5051.085 746.970 5051.685 ;
        RECT 748.000 5051.085 1213.000 5051.685 ;
        RECT 1213.965 5051.085 1291.970 5051.685 ;
        RECT 1293.000 5051.085 1758.000 5051.685 ;
        RECT 1758.965 5051.085 1836.970 5051.685 ;
        RECT 1838.000 5051.085 2303.000 5051.685 ;
        RECT 2303.965 5051.085 2381.970 5051.685 ;
        RECT 2383.000 5051.085 2848.000 5051.685 ;
        RECT 2848.965 5051.085 2922.035 5051.685 ;
        RECT 2923.000 5051.085 3588.000 5051.685 ;
        RECT 0.000 5045.835 202.330 5051.085 ;
      LAYER met4 ;
        RECT 202.730 5046.235 669.270 5050.685 ;
      LAYER met4 ;
        RECT 669.670 5045.835 746.330 5051.085 ;
      LAYER met4 ;
        RECT 746.730 5046.235 1214.270 5050.685 ;
      LAYER met4 ;
        RECT 1214.670 5045.835 1291.330 5051.085 ;
      LAYER met4 ;
        RECT 1291.730 5046.235 1759.270 5050.685 ;
      LAYER met4 ;
        RECT 1759.670 5045.835 1836.330 5051.085 ;
      LAYER met4 ;
        RECT 1836.730 5046.235 2304.270 5050.685 ;
      LAYER met4 ;
        RECT 2304.670 5045.835 2381.330 5051.085 ;
      LAYER met4 ;
        RECT 2381.730 5046.235 2849.270 5050.685 ;
      LAYER met4 ;
        RECT 2849.670 5045.835 2921.330 5051.085 ;
      LAYER met4 ;
        RECT 2921.730 5046.235 3389.625 5050.685 ;
      LAYER met4 ;
        RECT 3390.025 5045.835 3588.000 5051.085 ;
        RECT 0.000 5045.135 202.745 5045.835 ;
        RECT 204.000 5045.135 668.000 5045.835 ;
        RECT 668.965 5045.135 746.970 5045.835 ;
        RECT 748.000 5045.135 1213.000 5045.835 ;
        RECT 1213.965 5045.135 1291.970 5045.835 ;
        RECT 1293.000 5045.135 1758.000 5045.835 ;
        RECT 1758.965 5045.135 1836.970 5045.835 ;
        RECT 1838.000 5045.135 2303.000 5045.835 ;
        RECT 2303.965 5045.135 2381.970 5045.835 ;
        RECT 2383.000 5045.135 2848.000 5045.835 ;
        RECT 2848.965 5045.135 2922.035 5045.835 ;
        RECT 2923.000 5045.135 3588.000 5045.835 ;
        RECT 0.000 5044.005 176.425 5045.135 ;
      LAYER met4 ;
        RECT 176.825 5044.405 670.610 5044.735 ;
      LAYER met4 ;
        RECT 671.010 5044.505 714.690 5045.135 ;
        RECT 0.000 5040.725 176.690 5044.005 ;
      LAYER met4 ;
        RECT 177.090 5041.125 704.440 5044.105 ;
      LAYER met4 ;
        RECT 0.000 5039.245 182.045 5040.725 ;
      LAYER met4 ;
        RECT 182.445 5039.645 204.000 5040.825 ;
      LAYER met4 ;
        RECT 204.000 5039.745 668.000 5040.725 ;
      LAYER met4 ;
        RECT 668.000 5039.645 669.270 5040.825 ;
      LAYER met4 ;
        RECT 704.840 5040.725 706.360 5044.505 ;
      LAYER met4 ;
        RECT 715.090 5044.405 1215.610 5044.735 ;
      LAYER met4 ;
        RECT 1216.010 5044.505 1259.690 5045.135 ;
      LAYER met4 ;
        RECT 706.760 5041.125 1249.440 5044.105 ;
      LAYER met4 ;
        RECT 669.670 5039.745 746.330 5040.725 ;
        RECT 0.000 5036.465 182.725 5039.245 ;
        RECT 0.000 5035.335 180.025 5036.465 ;
      LAYER met4 ;
        RECT 183.125 5036.365 720.145 5039.345 ;
      LAYER met4 ;
        RECT 720.545 5036.465 722.065 5039.745 ;
      LAYER met4 ;
        RECT 746.730 5039.645 748.000 5040.825 ;
      LAYER met4 ;
        RECT 748.000 5039.745 1213.000 5040.725 ;
      LAYER met4 ;
        RECT 1213.000 5039.645 1214.270 5040.825 ;
      LAYER met4 ;
        RECT 1249.840 5040.725 1251.360 5044.505 ;
      LAYER met4 ;
        RECT 1260.090 5044.405 1760.610 5044.735 ;
      LAYER met4 ;
        RECT 1761.010 5044.505 1804.690 5045.135 ;
      LAYER met4 ;
        RECT 1251.760 5041.125 1794.440 5044.105 ;
      LAYER met4 ;
        RECT 1214.670 5039.745 1291.330 5040.725 ;
      LAYER met4 ;
        RECT 722.465 5036.365 1265.145 5039.345 ;
      LAYER met4 ;
        RECT 1265.545 5036.465 1267.065 5039.745 ;
      LAYER met4 ;
        RECT 1291.730 5039.645 1293.000 5040.825 ;
      LAYER met4 ;
        RECT 1293.000 5039.745 1758.000 5040.725 ;
      LAYER met4 ;
        RECT 1758.000 5039.645 1759.270 5040.825 ;
      LAYER met4 ;
        RECT 1794.840 5040.725 1796.360 5044.505 ;
      LAYER met4 ;
        RECT 1805.090 5044.405 2305.610 5044.735 ;
      LAYER met4 ;
        RECT 2306.010 5044.505 2349.690 5045.135 ;
      LAYER met4 ;
        RECT 1796.760 5041.125 2339.440 5044.105 ;
      LAYER met4 ;
        RECT 1759.670 5039.745 1836.330 5040.725 ;
      LAYER met4 ;
        RECT 1267.465 5036.365 1810.145 5039.345 ;
      LAYER met4 ;
        RECT 1810.545 5036.465 1812.065 5039.745 ;
      LAYER met4 ;
        RECT 1836.730 5039.645 1838.000 5040.825 ;
      LAYER met4 ;
        RECT 1838.000 5039.745 2303.000 5040.725 ;
      LAYER met4 ;
        RECT 2303.000 5039.645 2304.270 5040.825 ;
      LAYER met4 ;
        RECT 2339.840 5040.725 2341.360 5044.505 ;
      LAYER met4 ;
        RECT 2350.090 5044.405 3411.175 5044.735 ;
        RECT 2341.760 5041.125 3410.910 5044.105 ;
      LAYER met4 ;
        RECT 3411.575 5044.005 3588.000 5045.135 ;
        RECT 2304.670 5039.745 2381.330 5040.725 ;
      LAYER met4 ;
        RECT 1812.465 5036.365 2355.145 5039.345 ;
      LAYER met4 ;
        RECT 2355.545 5036.465 2357.065 5039.745 ;
      LAYER met4 ;
        RECT 2381.730 5039.645 2383.000 5040.825 ;
      LAYER met4 ;
        RECT 2383.000 5039.745 2848.000 5040.725 ;
      LAYER met4 ;
        RECT 2848.000 5039.645 2849.270 5040.825 ;
      LAYER met4 ;
        RECT 2849.670 5039.745 2921.330 5040.725 ;
      LAYER met4 ;
        RECT 2921.730 5039.645 2923.000 5040.825 ;
      LAYER met4 ;
        RECT 2923.000 5039.745 3388.000 5040.725 ;
      LAYER met4 ;
        RECT 3388.000 5039.645 3409.550 5040.825 ;
      LAYER met4 ;
        RECT 3411.310 5040.725 3588.000 5044.005 ;
      LAYER met4 ;
        RECT 2357.465 5036.365 3408.935 5039.345 ;
      LAYER met4 ;
        RECT 3409.950 5039.245 3588.000 5040.725 ;
      LAYER met4 ;
        RECT 180.425 5035.735 670.610 5036.065 ;
      LAYER met4 ;
        RECT 671.010 5035.335 714.690 5035.965 ;
      LAYER met4 ;
        RECT 715.090 5035.735 1215.610 5036.065 ;
      LAYER met4 ;
        RECT 1216.010 5035.335 1259.690 5035.965 ;
      LAYER met4 ;
        RECT 1260.090 5035.735 1760.610 5036.065 ;
      LAYER met4 ;
        RECT 1761.010 5035.335 1804.690 5035.965 ;
      LAYER met4 ;
        RECT 1805.090 5035.735 2305.610 5036.065 ;
      LAYER met4 ;
        RECT 2306.010 5035.335 2349.690 5035.965 ;
      LAYER met4 ;
        RECT 2350.090 5035.735 3407.575 5036.065 ;
      LAYER met4 ;
        RECT 3409.335 5035.965 3588.000 5039.245 ;
        RECT 3407.975 5035.335 3588.000 5035.965 ;
        RECT 0.000 5034.635 202.745 5035.335 ;
        RECT 668.965 5034.635 746.970 5035.335 ;
        RECT 1213.965 5034.635 1291.970 5035.335 ;
        RECT 1758.965 5034.635 1836.970 5035.335 ;
        RECT 2303.965 5034.635 2381.970 5035.335 ;
        RECT 2848.965 5034.635 2922.035 5035.335 ;
        RECT 3388.000 5034.635 3588.000 5035.335 ;
        RECT 0.000 5029.185 202.330 5034.635 ;
      LAYER met4 ;
        RECT 202.730 5029.585 669.270 5034.235 ;
      LAYER met4 ;
        RECT 669.670 5029.185 746.330 5034.635 ;
      LAYER met4 ;
        RECT 746.730 5029.585 1214.270 5034.235 ;
      LAYER met4 ;
        RECT 1214.670 5029.185 1291.330 5034.635 ;
      LAYER met4 ;
        RECT 1291.730 5029.585 1759.270 5034.235 ;
      LAYER met4 ;
        RECT 1759.670 5029.185 1836.330 5034.635 ;
      LAYER met4 ;
        RECT 1836.730 5029.585 2304.270 5034.235 ;
      LAYER met4 ;
        RECT 2304.670 5029.185 2381.330 5034.635 ;
      LAYER met4 ;
        RECT 2381.730 5029.585 2849.270 5034.235 ;
      LAYER met4 ;
        RECT 2849.670 5029.185 2921.330 5034.635 ;
      LAYER met4 ;
        RECT 2921.730 5029.585 3389.475 5034.235 ;
      LAYER met4 ;
        RECT 3389.875 5029.185 3588.000 5034.635 ;
        RECT 0.000 5028.585 202.745 5029.185 ;
        RECT 668.965 5028.585 746.970 5029.185 ;
        RECT 1213.965 5028.585 1291.970 5029.185 ;
        RECT 1758.965 5028.585 1836.970 5029.185 ;
        RECT 2303.965 5028.585 2381.970 5029.185 ;
        RECT 2848.965 5028.585 2922.035 5029.185 ;
        RECT 3388.000 5028.585 3588.000 5029.185 ;
        RECT 0.000 5024.335 202.330 5028.585 ;
      LAYER met4 ;
        RECT 202.730 5024.735 669.270 5028.185 ;
      LAYER met4 ;
        RECT 669.670 5024.335 746.330 5028.585 ;
      LAYER met4 ;
        RECT 746.730 5024.735 1214.270 5028.185 ;
      LAYER met4 ;
        RECT 1214.670 5024.335 1291.330 5028.585 ;
      LAYER met4 ;
        RECT 1291.730 5024.735 1759.270 5028.185 ;
      LAYER met4 ;
        RECT 1759.670 5024.335 1836.330 5028.585 ;
      LAYER met4 ;
        RECT 1836.730 5024.735 2304.270 5028.185 ;
      LAYER met4 ;
        RECT 2304.670 5024.335 2381.330 5028.585 ;
      LAYER met4 ;
        RECT 2381.730 5024.735 2849.270 5028.185 ;
      LAYER met4 ;
        RECT 2849.670 5024.335 2921.330 5028.585 ;
      LAYER met4 ;
        RECT 2921.730 5024.735 3389.335 5028.185 ;
      LAYER met4 ;
        RECT 3389.735 5024.335 3588.000 5028.585 ;
        RECT 0.000 5023.735 202.745 5024.335 ;
        RECT 668.965 5023.735 746.970 5024.335 ;
        RECT 1213.965 5023.735 1291.970 5024.335 ;
        RECT 1758.965 5023.735 1836.970 5024.335 ;
        RECT 2303.965 5023.735 2381.970 5024.335 ;
        RECT 2848.965 5023.735 2922.035 5024.335 ;
        RECT 3388.000 5023.735 3588.000 5024.335 ;
        RECT 0.000 5019.485 202.330 5023.735 ;
      LAYER met4 ;
        RECT 202.730 5019.885 669.270 5023.335 ;
      LAYER met4 ;
        RECT 669.670 5019.485 746.330 5023.735 ;
      LAYER met4 ;
        RECT 746.730 5019.885 1214.270 5023.335 ;
      LAYER met4 ;
        RECT 1214.670 5019.485 1291.330 5023.735 ;
      LAYER met4 ;
        RECT 1291.730 5019.885 1759.270 5023.335 ;
      LAYER met4 ;
        RECT 1759.670 5019.485 1836.330 5023.735 ;
      LAYER met4 ;
        RECT 1836.730 5019.885 2304.270 5023.335 ;
      LAYER met4 ;
        RECT 2304.670 5019.485 2381.330 5023.735 ;
      LAYER met4 ;
        RECT 2381.730 5019.885 2849.270 5023.335 ;
      LAYER met4 ;
        RECT 2849.670 5019.485 2921.330 5023.735 ;
      LAYER met4 ;
        RECT 2921.730 5019.885 3389.385 5023.335 ;
      LAYER met4 ;
        RECT 3389.785 5019.485 3588.000 5023.735 ;
        RECT 0.000 5018.885 202.745 5019.485 ;
        RECT 668.965 5018.885 746.970 5019.485 ;
        RECT 1213.965 5018.885 1291.970 5019.485 ;
        RECT 1758.965 5018.885 1836.970 5019.485 ;
        RECT 2303.965 5018.885 2381.970 5019.485 ;
        RECT 2848.965 5018.885 2922.035 5019.485 ;
        RECT 3388.000 5018.885 3588.000 5019.485 ;
        RECT 0.000 5013.435 202.330 5018.885 ;
      LAYER met4 ;
        RECT 202.730 5013.835 669.270 5018.485 ;
      LAYER met4 ;
        RECT 669.670 5013.435 746.330 5018.885 ;
      LAYER met4 ;
        RECT 746.730 5013.835 1214.270 5018.485 ;
      LAYER met4 ;
        RECT 1214.670 5013.435 1291.330 5018.885 ;
      LAYER met4 ;
        RECT 1291.730 5013.835 1759.270 5018.485 ;
      LAYER met4 ;
        RECT 1759.670 5013.435 1836.330 5018.885 ;
      LAYER met4 ;
        RECT 1836.730 5013.835 2304.270 5018.485 ;
      LAYER met4 ;
        RECT 2304.670 5013.435 2381.330 5018.885 ;
      LAYER met4 ;
        RECT 2381.730 5013.835 2849.270 5018.485 ;
      LAYER met4 ;
        RECT 2849.670 5013.435 2921.330 5018.885 ;
      LAYER met4 ;
        RECT 2921.730 5013.835 3389.600 5018.485 ;
      LAYER met4 ;
        RECT 3390.000 5013.435 3588.000 5018.885 ;
        RECT 0.000 5012.835 202.745 5013.435 ;
        RECT 668.965 5012.835 746.970 5013.435 ;
        RECT 1213.965 5012.835 1291.970 5013.435 ;
        RECT 1758.965 5012.835 1836.970 5013.435 ;
        RECT 2303.965 5012.835 2381.970 5013.435 ;
        RECT 2848.965 5012.835 2922.035 5013.435 ;
        RECT 3388.000 5012.835 3588.000 5013.435 ;
        RECT 0.000 5011.575 202.330 5012.835 ;
        RECT 0.000 4991.045 142.865 5011.575 ;
        RECT 143.995 5011.310 202.330 5011.575 ;
        RECT 0.000 4989.835 104.600 4991.045 ;
      LAYER met4 ;
        RECT 0.000 4988.000 24.215 4989.435 ;
      LAYER met4 ;
        RECT 24.615 4988.000 104.600 4989.835 ;
        RECT 0.000 4459.000 25.965 4988.000 ;
        RECT 102.965 4983.000 105.000 4988.000 ;
      LAYER met4 ;
        RECT 105.000 4983.000 129.965 4990.645 ;
      LAYER met4 ;
        RECT 130.365 4990.025 142.865 4991.045 ;
        RECT 130.365 4989.880 136.915 4990.025 ;
        RECT 130.365 4988.000 131.065 4989.880 ;
        RECT 129.965 4983.000 131.065 4988.000 ;
        RECT 102.965 4980.000 131.065 4983.000 ;
        RECT 102.965 4978.000 105.000 4980.000 ;
      LAYER met4 ;
        RECT 105.000 4978.000 129.965 4980.000 ;
      LAYER met4 ;
        RECT 129.965 4978.000 131.065 4980.000 ;
        RECT 102.965 4960.000 131.065 4978.000 ;
        RECT 102.965 4958.000 105.000 4960.000 ;
      LAYER met4 ;
        RECT 105.000 4958.000 129.965 4960.000 ;
      LAYER met4 ;
        RECT 129.965 4958.000 131.065 4960.000 ;
        RECT 102.965 4940.000 131.065 4958.000 ;
        RECT 102.965 4938.000 105.000 4940.000 ;
      LAYER met4 ;
        RECT 105.000 4938.000 129.965 4940.000 ;
      LAYER met4 ;
        RECT 129.965 4938.000 131.065 4940.000 ;
        RECT 102.965 4920.000 131.065 4938.000 ;
        RECT 102.965 4918.000 105.000 4920.000 ;
      LAYER met4 ;
        RECT 105.000 4918.000 129.965 4920.000 ;
      LAYER met4 ;
        RECT 129.965 4918.000 131.065 4920.000 ;
        RECT 102.965 4900.000 131.065 4918.000 ;
        RECT 102.965 4898.000 105.000 4900.000 ;
      LAYER met4 ;
        RECT 105.000 4898.000 129.965 4900.000 ;
      LAYER met4 ;
        RECT 129.965 4898.000 131.065 4900.000 ;
        RECT 102.965 4880.000 131.065 4898.000 ;
        RECT 102.965 4878.000 105.000 4880.000 ;
      LAYER met4 ;
        RECT 105.000 4878.000 129.965 4880.000 ;
      LAYER met4 ;
        RECT 129.965 4878.000 131.065 4880.000 ;
        RECT 102.965 4860.000 131.065 4878.000 ;
        RECT 102.965 4858.000 105.000 4860.000 ;
      LAYER met4 ;
        RECT 105.000 4858.000 129.965 4860.000 ;
      LAYER met4 ;
        RECT 129.965 4858.000 131.065 4860.000 ;
        RECT 102.965 4840.000 131.065 4858.000 ;
        RECT 102.965 4838.000 105.000 4840.000 ;
      LAYER met4 ;
        RECT 105.000 4838.000 129.965 4840.000 ;
      LAYER met4 ;
        RECT 129.965 4838.000 131.065 4840.000 ;
        RECT 102.965 4820.000 131.065 4838.000 ;
        RECT 102.965 4818.000 105.000 4820.000 ;
      LAYER met4 ;
        RECT 105.000 4818.000 129.965 4820.000 ;
      LAYER met4 ;
        RECT 129.965 4818.000 131.065 4820.000 ;
        RECT 102.965 4800.000 131.065 4818.000 ;
        RECT 102.965 4798.000 105.000 4800.000 ;
      LAYER met4 ;
        RECT 105.000 4798.000 129.965 4800.000 ;
      LAYER met4 ;
        RECT 129.965 4798.000 131.065 4800.000 ;
        RECT 102.965 4780.000 131.065 4798.000 ;
        RECT 102.965 4778.000 105.000 4780.000 ;
      LAYER met4 ;
        RECT 105.000 4778.000 129.965 4780.000 ;
      LAYER met4 ;
        RECT 129.965 4778.000 131.065 4780.000 ;
        RECT 102.965 4760.000 131.065 4778.000 ;
        RECT 102.965 4758.000 105.000 4760.000 ;
      LAYER met4 ;
        RECT 105.000 4758.000 129.965 4760.000 ;
      LAYER met4 ;
        RECT 129.965 4758.000 131.065 4760.000 ;
        RECT 102.965 4740.000 131.065 4758.000 ;
        RECT 102.965 4738.000 105.000 4740.000 ;
      LAYER met4 ;
        RECT 105.000 4738.000 129.965 4740.000 ;
      LAYER met4 ;
        RECT 129.965 4738.000 131.065 4740.000 ;
        RECT 102.965 4720.000 131.065 4738.000 ;
        RECT 102.965 4718.000 105.000 4720.000 ;
      LAYER met4 ;
        RECT 105.000 4718.000 129.965 4720.000 ;
      LAYER met4 ;
        RECT 129.965 4718.000 131.065 4720.000 ;
        RECT 102.965 4700.000 131.065 4718.000 ;
        RECT 102.965 4698.000 105.000 4700.000 ;
      LAYER met4 ;
        RECT 105.000 4698.000 129.965 4700.000 ;
      LAYER met4 ;
        RECT 129.965 4698.000 131.065 4700.000 ;
        RECT 102.965 4680.000 131.065 4698.000 ;
        RECT 102.965 4678.000 105.000 4680.000 ;
      LAYER met4 ;
        RECT 105.000 4678.000 129.965 4680.000 ;
      LAYER met4 ;
        RECT 129.965 4678.000 131.065 4680.000 ;
        RECT 102.965 4660.000 131.065 4678.000 ;
        RECT 102.965 4658.000 105.000 4660.000 ;
      LAYER met4 ;
        RECT 105.000 4658.000 129.965 4660.000 ;
      LAYER met4 ;
        RECT 129.965 4658.000 131.065 4660.000 ;
        RECT 102.965 4640.000 131.065 4658.000 ;
        RECT 102.965 4638.000 105.000 4640.000 ;
      LAYER met4 ;
        RECT 105.000 4638.000 129.965 4640.000 ;
      LAYER met4 ;
        RECT 129.965 4638.000 131.065 4640.000 ;
        RECT 102.965 4620.000 131.065 4638.000 ;
        RECT 102.965 4618.000 105.000 4620.000 ;
      LAYER met4 ;
        RECT 105.000 4618.000 129.965 4620.000 ;
      LAYER met4 ;
        RECT 129.965 4618.000 131.065 4620.000 ;
        RECT 102.965 4600.000 131.065 4618.000 ;
        RECT 102.965 4598.000 105.000 4600.000 ;
      LAYER met4 ;
        RECT 105.000 4598.000 129.965 4600.000 ;
      LAYER met4 ;
        RECT 129.965 4598.000 131.065 4600.000 ;
        RECT 102.965 4580.000 131.065 4598.000 ;
        RECT 102.965 4578.000 105.000 4580.000 ;
      LAYER met4 ;
        RECT 105.000 4578.000 129.965 4580.000 ;
      LAYER met4 ;
        RECT 129.965 4578.000 131.065 4580.000 ;
        RECT 102.965 4560.000 131.065 4578.000 ;
        RECT 102.965 4558.000 105.000 4560.000 ;
      LAYER met4 ;
        RECT 105.000 4558.000 129.965 4560.000 ;
      LAYER met4 ;
        RECT 129.965 4558.000 131.065 4560.000 ;
        RECT 102.965 4540.000 131.065 4558.000 ;
        RECT 102.965 4538.000 105.000 4540.000 ;
      LAYER met4 ;
        RECT 105.000 4538.000 129.965 4540.000 ;
      LAYER met4 ;
        RECT 129.965 4538.000 131.065 4540.000 ;
        RECT 102.965 4520.000 131.065 4538.000 ;
        RECT 102.965 4518.000 105.000 4520.000 ;
      LAYER met4 ;
        RECT 105.000 4518.000 129.965 4520.000 ;
      LAYER met4 ;
        RECT 129.965 4518.000 131.065 4520.000 ;
        RECT 102.965 4500.000 131.065 4518.000 ;
        RECT 102.965 4498.000 105.000 4500.000 ;
      LAYER met4 ;
        RECT 105.000 4498.000 129.965 4500.000 ;
      LAYER met4 ;
        RECT 129.965 4498.000 131.065 4500.000 ;
        RECT 102.965 4480.000 131.065 4498.000 ;
        RECT 102.965 4478.000 105.000 4480.000 ;
      LAYER met4 ;
        RECT 105.000 4478.000 129.965 4480.000 ;
      LAYER met4 ;
        RECT 129.965 4478.000 131.065 4480.000 ;
        RECT 102.965 4460.000 131.065 4478.000 ;
        RECT 102.965 4459.000 105.000 4460.000 ;
      LAYER met4 ;
        RECT 0.000 4457.730 24.215 4459.000 ;
      LAYER met4 ;
        RECT 24.615 4457.330 104.600 4458.035 ;
      LAYER met4 ;
        RECT 105.000 4457.730 129.965 4460.000 ;
      LAYER met4 ;
        RECT 129.965 4459.000 131.065 4460.000 ;
        RECT 130.365 4457.330 131.065 4458.035 ;
      LAYER met4 ;
        RECT 131.465 4457.730 135.915 4989.480 ;
      LAYER met4 ;
        RECT 136.315 4988.000 136.915 4989.880 ;
        RECT 136.315 4459.000 136.915 4984.000 ;
        RECT 136.315 4457.330 136.915 4458.035 ;
      LAYER met4 ;
        RECT 137.315 4457.730 141.765 4989.625 ;
      LAYER met4 ;
        RECT 142.165 4459.000 142.865 4990.025 ;
        RECT 142.165 4457.330 142.865 4458.035 ;
        RECT 0.000 4385.670 142.865 4457.330 ;
      LAYER met4 ;
        RECT 0.000 4384.000 24.215 4385.270 ;
      LAYER met4 ;
        RECT 24.615 4384.965 104.600 4385.670 ;
        RECT 0.000 3855.000 25.965 4384.000 ;
        RECT 102.965 4379.000 105.000 4384.000 ;
      LAYER met4 ;
        RECT 105.000 4379.000 129.965 4385.270 ;
      LAYER met4 ;
        RECT 130.365 4384.965 131.065 4385.670 ;
        RECT 129.965 4379.000 131.065 4384.000 ;
        RECT 102.965 4376.000 131.065 4379.000 ;
        RECT 102.965 4374.000 105.000 4376.000 ;
      LAYER met4 ;
        RECT 105.000 4374.000 129.965 4376.000 ;
      LAYER met4 ;
        RECT 129.965 4374.000 131.065 4376.000 ;
        RECT 102.965 4356.000 131.065 4374.000 ;
        RECT 102.965 4354.000 105.000 4356.000 ;
      LAYER met4 ;
        RECT 105.000 4354.000 129.965 4356.000 ;
      LAYER met4 ;
        RECT 129.965 4354.000 131.065 4356.000 ;
        RECT 102.965 4336.000 131.065 4354.000 ;
        RECT 102.965 4334.000 105.000 4336.000 ;
      LAYER met4 ;
        RECT 105.000 4334.000 129.965 4336.000 ;
      LAYER met4 ;
        RECT 129.965 4334.000 131.065 4336.000 ;
        RECT 102.965 4316.000 131.065 4334.000 ;
        RECT 102.965 4314.000 105.000 4316.000 ;
      LAYER met4 ;
        RECT 105.000 4314.000 129.965 4316.000 ;
      LAYER met4 ;
        RECT 129.965 4314.000 131.065 4316.000 ;
        RECT 102.965 4296.000 131.065 4314.000 ;
        RECT 102.965 4294.000 105.000 4296.000 ;
      LAYER met4 ;
        RECT 105.000 4294.000 129.965 4296.000 ;
      LAYER met4 ;
        RECT 129.965 4294.000 131.065 4296.000 ;
        RECT 102.965 4276.000 131.065 4294.000 ;
        RECT 102.965 4274.000 105.000 4276.000 ;
      LAYER met4 ;
        RECT 105.000 4274.000 129.965 4276.000 ;
      LAYER met4 ;
        RECT 129.965 4274.000 131.065 4276.000 ;
        RECT 102.965 4256.000 131.065 4274.000 ;
        RECT 102.965 4254.000 105.000 4256.000 ;
      LAYER met4 ;
        RECT 105.000 4254.000 129.965 4256.000 ;
      LAYER met4 ;
        RECT 129.965 4254.000 131.065 4256.000 ;
        RECT 102.965 4236.000 131.065 4254.000 ;
        RECT 102.965 4234.000 105.000 4236.000 ;
      LAYER met4 ;
        RECT 105.000 4234.000 129.965 4236.000 ;
      LAYER met4 ;
        RECT 129.965 4234.000 131.065 4236.000 ;
        RECT 102.965 4216.000 131.065 4234.000 ;
        RECT 102.965 4214.000 105.000 4216.000 ;
      LAYER met4 ;
        RECT 105.000 4214.000 129.965 4216.000 ;
      LAYER met4 ;
        RECT 129.965 4214.000 131.065 4216.000 ;
        RECT 102.965 4196.000 131.065 4214.000 ;
        RECT 102.965 4194.000 105.000 4196.000 ;
      LAYER met4 ;
        RECT 105.000 4194.000 129.965 4196.000 ;
      LAYER met4 ;
        RECT 129.965 4194.000 131.065 4196.000 ;
        RECT 102.965 4176.000 131.065 4194.000 ;
        RECT 102.965 4174.000 105.000 4176.000 ;
      LAYER met4 ;
        RECT 105.000 4174.000 129.965 4176.000 ;
      LAYER met4 ;
        RECT 129.965 4174.000 131.065 4176.000 ;
        RECT 102.965 4156.000 131.065 4174.000 ;
        RECT 102.965 4154.000 105.000 4156.000 ;
      LAYER met4 ;
        RECT 105.000 4154.000 129.965 4156.000 ;
      LAYER met4 ;
        RECT 129.965 4154.000 131.065 4156.000 ;
        RECT 102.965 4136.000 131.065 4154.000 ;
        RECT 102.965 4134.000 105.000 4136.000 ;
      LAYER met4 ;
        RECT 105.000 4134.000 129.965 4136.000 ;
      LAYER met4 ;
        RECT 129.965 4134.000 131.065 4136.000 ;
        RECT 102.965 4116.000 131.065 4134.000 ;
        RECT 102.965 4114.000 105.000 4116.000 ;
      LAYER met4 ;
        RECT 105.000 4114.000 129.965 4116.000 ;
      LAYER met4 ;
        RECT 129.965 4114.000 131.065 4116.000 ;
        RECT 102.965 4096.000 131.065 4114.000 ;
        RECT 102.965 4094.000 105.000 4096.000 ;
      LAYER met4 ;
        RECT 105.000 4094.000 129.965 4096.000 ;
      LAYER met4 ;
        RECT 129.965 4094.000 131.065 4096.000 ;
        RECT 102.965 4076.000 131.065 4094.000 ;
        RECT 102.965 4074.000 105.000 4076.000 ;
      LAYER met4 ;
        RECT 105.000 4074.000 129.965 4076.000 ;
      LAYER met4 ;
        RECT 129.965 4074.000 131.065 4076.000 ;
        RECT 102.965 4056.000 131.065 4074.000 ;
        RECT 102.965 4054.000 105.000 4056.000 ;
      LAYER met4 ;
        RECT 105.000 4054.000 129.965 4056.000 ;
      LAYER met4 ;
        RECT 129.965 4054.000 131.065 4056.000 ;
        RECT 102.965 4036.000 131.065 4054.000 ;
        RECT 102.965 4034.000 105.000 4036.000 ;
      LAYER met4 ;
        RECT 105.000 4034.000 129.965 4036.000 ;
      LAYER met4 ;
        RECT 129.965 4034.000 131.065 4036.000 ;
        RECT 102.965 4016.000 131.065 4034.000 ;
        RECT 102.965 4014.000 105.000 4016.000 ;
      LAYER met4 ;
        RECT 105.000 4014.000 129.965 4016.000 ;
      LAYER met4 ;
        RECT 129.965 4014.000 131.065 4016.000 ;
        RECT 102.965 3996.000 131.065 4014.000 ;
        RECT 102.965 3994.000 105.000 3996.000 ;
      LAYER met4 ;
        RECT 105.000 3994.000 129.965 3996.000 ;
      LAYER met4 ;
        RECT 129.965 3994.000 131.065 3996.000 ;
        RECT 102.965 3976.000 131.065 3994.000 ;
        RECT 102.965 3974.000 105.000 3976.000 ;
      LAYER met4 ;
        RECT 105.000 3974.000 129.965 3976.000 ;
      LAYER met4 ;
        RECT 129.965 3974.000 131.065 3976.000 ;
        RECT 102.965 3956.000 131.065 3974.000 ;
        RECT 102.965 3954.000 105.000 3956.000 ;
      LAYER met4 ;
        RECT 105.000 3954.000 129.965 3956.000 ;
      LAYER met4 ;
        RECT 129.965 3954.000 131.065 3956.000 ;
        RECT 102.965 3936.000 131.065 3954.000 ;
        RECT 102.965 3934.000 105.000 3936.000 ;
      LAYER met4 ;
        RECT 105.000 3934.000 129.965 3936.000 ;
      LAYER met4 ;
        RECT 129.965 3934.000 131.065 3936.000 ;
        RECT 102.965 3916.000 131.065 3934.000 ;
        RECT 102.965 3914.000 105.000 3916.000 ;
      LAYER met4 ;
        RECT 105.000 3914.000 129.965 3916.000 ;
      LAYER met4 ;
        RECT 129.965 3914.000 131.065 3916.000 ;
        RECT 102.965 3896.000 131.065 3914.000 ;
        RECT 102.965 3894.000 105.000 3896.000 ;
      LAYER met4 ;
        RECT 105.000 3894.000 129.965 3896.000 ;
      LAYER met4 ;
        RECT 129.965 3894.000 131.065 3896.000 ;
        RECT 102.965 3876.000 131.065 3894.000 ;
        RECT 102.965 3874.000 105.000 3876.000 ;
      LAYER met4 ;
        RECT 105.000 3874.000 129.965 3876.000 ;
      LAYER met4 ;
        RECT 129.965 3874.000 131.065 3876.000 ;
        RECT 102.965 3856.000 131.065 3874.000 ;
        RECT 102.965 3855.000 105.000 3856.000 ;
      LAYER met4 ;
        RECT 0.000 3853.730 24.215 3855.000 ;
      LAYER met4 ;
        RECT 24.615 3853.330 104.600 3853.970 ;
      LAYER met4 ;
        RECT 105.000 3853.730 129.965 3856.000 ;
      LAYER met4 ;
        RECT 129.965 3855.000 131.065 3856.000 ;
        RECT 130.365 3853.330 131.065 3853.970 ;
      LAYER met4 ;
        RECT 131.465 3853.730 135.915 4385.270 ;
      LAYER met4 ;
        RECT 136.315 4384.965 136.915 4385.670 ;
        RECT 136.315 3855.000 136.915 4380.000 ;
        RECT 136.315 3853.330 136.915 3853.970 ;
      LAYER met4 ;
        RECT 137.315 3853.730 141.765 4385.270 ;
      LAYER met4 ;
        RECT 142.165 4384.965 142.865 4385.670 ;
        RECT 142.165 3855.000 142.865 4384.000 ;
        RECT 142.165 3853.330 142.865 3853.970 ;
        RECT 0.000 3821.690 142.865 3853.330 ;
      LAYER met4 ;
        RECT 143.265 3822.090 143.595 5011.175 ;
      LAYER met4 ;
        RECT 0.000 3813.360 143.495 3821.690 ;
      LAYER met4 ;
        RECT 143.895 3813.760 146.875 5010.910 ;
      LAYER met4 ;
        RECT 147.275 5009.950 202.330 5011.310 ;
      LAYER met4 ;
        RECT 147.175 4988.000 148.355 5009.550 ;
      LAYER met4 ;
        RECT 148.755 5009.335 202.330 5009.950 ;
        RECT 147.275 4459.000 148.255 4988.000 ;
      LAYER met4 ;
        RECT 147.175 4457.730 148.355 4459.000 ;
      LAYER met4 ;
        RECT 147.275 4385.670 148.255 4457.330 ;
      LAYER met4 ;
        RECT 147.175 4384.000 148.355 4385.270 ;
      LAYER met4 ;
        RECT 147.275 3855.000 148.255 4384.000 ;
      LAYER met4 ;
        RECT 147.175 3853.730 148.355 3855.000 ;
      LAYER met4 ;
        RECT 147.275 3829.065 148.255 3853.330 ;
      LAYER met4 ;
        RECT 148.655 3829.465 151.635 5008.935 ;
      LAYER met4 ;
        RECT 152.035 5007.975 202.330 5009.335 ;
        RECT 147.275 3827.545 151.535 3829.065 ;
        RECT 147.275 3813.360 148.255 3827.545 ;
        RECT 0.000 3811.840 148.255 3813.360 ;
        RECT 0.000 3778.010 143.495 3811.840 ;
        RECT 0.000 3776.670 142.865 3778.010 ;
      LAYER met4 ;
        RECT 0.000 3775.000 24.215 3776.270 ;
      LAYER met4 ;
        RECT 24.615 3775.965 104.600 3776.670 ;
        RECT 0.000 3247.000 25.965 3775.000 ;
        RECT 102.965 3771.000 105.000 3775.000 ;
      LAYER met4 ;
        RECT 105.000 3771.000 129.965 3776.270 ;
      LAYER met4 ;
        RECT 130.365 3775.965 131.065 3776.670 ;
        RECT 129.965 3771.000 131.065 3775.000 ;
        RECT 102.965 3768.000 131.065 3771.000 ;
        RECT 102.965 3766.000 105.000 3768.000 ;
      LAYER met4 ;
        RECT 105.000 3766.000 129.965 3768.000 ;
      LAYER met4 ;
        RECT 129.965 3766.000 131.065 3768.000 ;
        RECT 102.965 3748.000 131.065 3766.000 ;
        RECT 102.965 3746.000 105.000 3748.000 ;
      LAYER met4 ;
        RECT 105.000 3746.000 129.965 3748.000 ;
      LAYER met4 ;
        RECT 129.965 3746.000 131.065 3748.000 ;
        RECT 102.965 3728.000 131.065 3746.000 ;
        RECT 102.965 3726.000 105.000 3728.000 ;
      LAYER met4 ;
        RECT 105.000 3726.000 129.965 3728.000 ;
      LAYER met4 ;
        RECT 129.965 3726.000 131.065 3728.000 ;
        RECT 102.965 3708.000 131.065 3726.000 ;
        RECT 102.965 3706.000 105.000 3708.000 ;
      LAYER met4 ;
        RECT 105.000 3706.000 129.965 3708.000 ;
      LAYER met4 ;
        RECT 129.965 3706.000 131.065 3708.000 ;
        RECT 102.965 3688.000 131.065 3706.000 ;
        RECT 102.965 3686.000 105.000 3688.000 ;
      LAYER met4 ;
        RECT 105.000 3686.000 129.965 3688.000 ;
      LAYER met4 ;
        RECT 129.965 3686.000 131.065 3688.000 ;
        RECT 102.965 3668.000 131.065 3686.000 ;
        RECT 102.965 3666.000 105.000 3668.000 ;
      LAYER met4 ;
        RECT 105.000 3666.000 129.965 3668.000 ;
      LAYER met4 ;
        RECT 129.965 3666.000 131.065 3668.000 ;
        RECT 102.965 3648.000 131.065 3666.000 ;
        RECT 102.965 3646.000 105.000 3648.000 ;
      LAYER met4 ;
        RECT 105.000 3646.000 129.965 3648.000 ;
      LAYER met4 ;
        RECT 129.965 3646.000 131.065 3648.000 ;
        RECT 102.965 3628.000 131.065 3646.000 ;
        RECT 102.965 3626.000 105.000 3628.000 ;
      LAYER met4 ;
        RECT 105.000 3626.000 129.965 3628.000 ;
      LAYER met4 ;
        RECT 129.965 3626.000 131.065 3628.000 ;
        RECT 102.965 3608.000 131.065 3626.000 ;
        RECT 102.965 3606.000 105.000 3608.000 ;
      LAYER met4 ;
        RECT 105.000 3606.000 129.965 3608.000 ;
      LAYER met4 ;
        RECT 129.965 3606.000 131.065 3608.000 ;
        RECT 102.965 3588.000 131.065 3606.000 ;
        RECT 102.965 3586.000 105.000 3588.000 ;
      LAYER met4 ;
        RECT 105.000 3586.000 129.965 3588.000 ;
      LAYER met4 ;
        RECT 129.965 3586.000 131.065 3588.000 ;
        RECT 102.965 3568.000 131.065 3586.000 ;
        RECT 102.965 3566.000 105.000 3568.000 ;
      LAYER met4 ;
        RECT 105.000 3566.000 129.965 3568.000 ;
      LAYER met4 ;
        RECT 129.965 3566.000 131.065 3568.000 ;
        RECT 102.965 3548.000 131.065 3566.000 ;
        RECT 102.965 3546.000 105.000 3548.000 ;
      LAYER met4 ;
        RECT 105.000 3546.000 129.965 3548.000 ;
      LAYER met4 ;
        RECT 129.965 3546.000 131.065 3548.000 ;
        RECT 102.965 3528.000 131.065 3546.000 ;
        RECT 102.965 3526.000 105.000 3528.000 ;
      LAYER met4 ;
        RECT 105.000 3526.000 129.965 3528.000 ;
      LAYER met4 ;
        RECT 129.965 3526.000 131.065 3528.000 ;
        RECT 102.965 3508.000 131.065 3526.000 ;
        RECT 102.965 3506.000 105.000 3508.000 ;
      LAYER met4 ;
        RECT 105.000 3506.000 129.965 3508.000 ;
      LAYER met4 ;
        RECT 129.965 3506.000 131.065 3508.000 ;
        RECT 102.965 3488.000 131.065 3506.000 ;
        RECT 102.965 3486.000 105.000 3488.000 ;
      LAYER met4 ;
        RECT 105.000 3486.000 129.965 3488.000 ;
      LAYER met4 ;
        RECT 129.965 3486.000 131.065 3488.000 ;
        RECT 102.965 3468.000 131.065 3486.000 ;
        RECT 102.965 3466.000 105.000 3468.000 ;
      LAYER met4 ;
        RECT 105.000 3466.000 129.965 3468.000 ;
      LAYER met4 ;
        RECT 129.965 3466.000 131.065 3468.000 ;
        RECT 102.965 3448.000 131.065 3466.000 ;
        RECT 102.965 3446.000 105.000 3448.000 ;
      LAYER met4 ;
        RECT 105.000 3446.000 129.965 3448.000 ;
      LAYER met4 ;
        RECT 129.965 3446.000 131.065 3448.000 ;
        RECT 102.965 3428.000 131.065 3446.000 ;
        RECT 102.965 3426.000 105.000 3428.000 ;
      LAYER met4 ;
        RECT 105.000 3426.000 129.965 3428.000 ;
      LAYER met4 ;
        RECT 129.965 3426.000 131.065 3428.000 ;
        RECT 102.965 3408.000 131.065 3426.000 ;
        RECT 102.965 3406.000 105.000 3408.000 ;
      LAYER met4 ;
        RECT 105.000 3406.000 129.965 3408.000 ;
      LAYER met4 ;
        RECT 129.965 3406.000 131.065 3408.000 ;
        RECT 102.965 3388.000 131.065 3406.000 ;
        RECT 102.965 3386.000 105.000 3388.000 ;
      LAYER met4 ;
        RECT 105.000 3386.000 129.965 3388.000 ;
      LAYER met4 ;
        RECT 129.965 3386.000 131.065 3388.000 ;
        RECT 102.965 3368.000 131.065 3386.000 ;
        RECT 102.965 3366.000 105.000 3368.000 ;
      LAYER met4 ;
        RECT 105.000 3366.000 129.965 3368.000 ;
      LAYER met4 ;
        RECT 129.965 3366.000 131.065 3368.000 ;
        RECT 102.965 3348.000 131.065 3366.000 ;
        RECT 102.965 3346.000 105.000 3348.000 ;
      LAYER met4 ;
        RECT 105.000 3346.000 129.965 3348.000 ;
      LAYER met4 ;
        RECT 129.965 3346.000 131.065 3348.000 ;
        RECT 102.965 3328.000 131.065 3346.000 ;
        RECT 102.965 3326.000 105.000 3328.000 ;
      LAYER met4 ;
        RECT 105.000 3326.000 129.965 3328.000 ;
      LAYER met4 ;
        RECT 129.965 3326.000 131.065 3328.000 ;
        RECT 102.965 3308.000 131.065 3326.000 ;
        RECT 102.965 3306.000 105.000 3308.000 ;
      LAYER met4 ;
        RECT 105.000 3306.000 129.965 3308.000 ;
      LAYER met4 ;
        RECT 129.965 3306.000 131.065 3308.000 ;
        RECT 102.965 3288.000 131.065 3306.000 ;
        RECT 102.965 3286.000 105.000 3288.000 ;
      LAYER met4 ;
        RECT 105.000 3286.000 129.965 3288.000 ;
      LAYER met4 ;
        RECT 129.965 3286.000 131.065 3288.000 ;
        RECT 102.965 3268.000 131.065 3286.000 ;
        RECT 102.965 3266.000 105.000 3268.000 ;
      LAYER met4 ;
        RECT 105.000 3266.000 129.965 3268.000 ;
      LAYER met4 ;
        RECT 129.965 3266.000 131.065 3268.000 ;
        RECT 102.965 3248.000 131.065 3266.000 ;
        RECT 102.965 3247.000 105.000 3248.000 ;
      LAYER met4 ;
        RECT 0.000 3245.730 24.215 3247.000 ;
      LAYER met4 ;
        RECT 24.615 3245.330 104.600 3245.970 ;
      LAYER met4 ;
        RECT 105.000 3245.730 129.965 3248.000 ;
      LAYER met4 ;
        RECT 129.965 3247.000 131.065 3248.000 ;
        RECT 130.365 3245.330 131.065 3245.970 ;
      LAYER met4 ;
        RECT 131.465 3245.730 135.915 3776.270 ;
      LAYER met4 ;
        RECT 136.315 3775.965 136.915 3776.670 ;
        RECT 136.315 3247.000 136.915 3772.000 ;
        RECT 136.315 3245.330 136.915 3245.970 ;
      LAYER met4 ;
        RECT 137.315 3245.730 141.765 3776.270 ;
      LAYER met4 ;
        RECT 142.165 3775.965 142.865 3776.670 ;
        RECT 142.165 3247.000 142.865 3775.000 ;
        RECT 142.165 3245.330 142.865 3245.970 ;
        RECT 0.000 3213.690 142.865 3245.330 ;
      LAYER met4 ;
        RECT 143.265 3214.090 143.595 3777.610 ;
      LAYER met4 ;
        RECT 0.000 3205.360 143.495 3213.690 ;
      LAYER met4 ;
        RECT 143.895 3205.760 146.875 3811.440 ;
      LAYER met4 ;
        RECT 147.275 3776.670 148.255 3811.840 ;
      LAYER met4 ;
        RECT 147.175 3775.000 148.355 3776.270 ;
      LAYER met4 ;
        RECT 147.275 3247.000 148.255 3775.000 ;
      LAYER met4 ;
        RECT 147.175 3245.730 148.355 3247.000 ;
      LAYER met4 ;
        RECT 147.275 3221.065 148.255 3245.330 ;
      LAYER met4 ;
        RECT 148.655 3221.465 151.635 3827.145 ;
        RECT 151.935 3822.090 152.265 5007.575 ;
      LAYER met4 ;
        RECT 152.665 5007.385 202.330 5007.975 ;
      LAYER met4 ;
        RECT 202.730 5007.785 669.270 5012.435 ;
      LAYER met4 ;
        RECT 669.670 5007.385 746.330 5012.835 ;
      LAYER met4 ;
        RECT 746.730 5007.785 1214.270 5012.435 ;
      LAYER met4 ;
        RECT 1214.670 5007.385 1291.330 5012.835 ;
      LAYER met4 ;
        RECT 1291.730 5007.785 1759.270 5012.435 ;
      LAYER met4 ;
        RECT 1759.670 5007.385 1836.330 5012.835 ;
      LAYER met4 ;
        RECT 1836.730 5007.785 2304.270 5012.435 ;
      LAYER met4 ;
        RECT 2304.670 5007.385 2381.330 5012.835 ;
      LAYER met4 ;
        RECT 2381.730 5007.785 2849.270 5012.435 ;
      LAYER met4 ;
        RECT 2849.670 5007.385 2921.330 5012.835 ;
      LAYER met4 ;
        RECT 2921.730 5007.785 3389.525 5012.435 ;
      LAYER met4 ;
        RECT 3389.925 5011.575 3588.000 5012.835 ;
        RECT 3389.925 5011.310 3444.005 5011.575 ;
        RECT 3389.925 5007.975 3440.725 5011.310 ;
        RECT 3389.925 5007.385 3435.335 5007.975 ;
        RECT 152.665 5006.785 202.745 5007.385 ;
        RECT 668.965 5006.785 746.970 5007.385 ;
        RECT 1213.965 5006.785 1291.970 5007.385 ;
        RECT 1758.965 5006.785 1836.970 5007.385 ;
        RECT 2303.965 5006.785 2381.970 5007.385 ;
        RECT 2848.965 5006.785 2922.035 5007.385 ;
        RECT 3388.000 5006.785 3435.335 5007.385 ;
        RECT 152.665 5002.535 202.345 5006.785 ;
      LAYER met4 ;
        RECT 202.745 5002.935 668.965 5006.385 ;
      LAYER met4 ;
        RECT 669.365 5002.535 746.570 5006.785 ;
      LAYER met4 ;
        RECT 746.970 5002.935 1213.965 5006.385 ;
      LAYER met4 ;
        RECT 1214.365 5002.535 1291.570 5006.785 ;
      LAYER met4 ;
        RECT 1291.970 5002.935 1758.965 5006.385 ;
      LAYER met4 ;
        RECT 1759.365 5002.535 1836.570 5006.785 ;
      LAYER met4 ;
        RECT 1836.970 5002.935 2303.965 5006.385 ;
      LAYER met4 ;
        RECT 2304.365 5002.535 2381.570 5006.785 ;
      LAYER met4 ;
        RECT 2381.970 5002.935 2848.965 5006.385 ;
      LAYER met4 ;
        RECT 2849.365 5002.535 2921.635 5006.785 ;
      LAYER met4 ;
        RECT 2922.035 5002.935 3389.470 5006.385 ;
      LAYER met4 ;
        RECT 3389.870 5002.535 3435.335 5006.785 ;
        RECT 152.665 5001.935 202.745 5002.535 ;
        RECT 668.965 5001.935 746.970 5002.535 ;
        RECT 1213.965 5001.935 1291.970 5002.535 ;
        RECT 1758.965 5001.935 1836.970 5002.535 ;
        RECT 2303.965 5001.935 2381.970 5002.535 ;
        RECT 2848.965 5001.935 2922.035 5002.535 ;
        RECT 3388.000 5001.935 3435.335 5002.535 ;
        RECT 152.665 4996.485 202.330 5001.935 ;
      LAYER met4 ;
        RECT 202.730 4996.885 669.270 5001.535 ;
      LAYER met4 ;
        RECT 669.670 4996.485 746.330 5001.935 ;
      LAYER met4 ;
        RECT 746.730 4996.885 1214.270 5001.535 ;
      LAYER met4 ;
        RECT 1214.670 4996.485 1291.330 5001.935 ;
      LAYER met4 ;
        RECT 1291.730 4996.885 1759.270 5001.535 ;
      LAYER met4 ;
        RECT 1759.670 4996.485 1836.330 5001.935 ;
      LAYER met4 ;
        RECT 1836.730 4996.885 2304.270 5001.535 ;
      LAYER met4 ;
        RECT 2304.670 4996.485 2381.330 5001.935 ;
      LAYER met4 ;
        RECT 2381.730 4996.885 2849.270 5001.535 ;
      LAYER met4 ;
        RECT 2849.670 4996.485 2921.330 5001.935 ;
      LAYER met4 ;
        RECT 2921.730 4996.885 3391.785 5001.535 ;
      LAYER met4 ;
        RECT 3392.185 4996.485 3435.335 5001.935 ;
        RECT 152.665 4995.885 202.745 4996.485 ;
        RECT 668.965 4995.885 746.970 4996.485 ;
        RECT 1213.965 4995.885 1291.970 4996.485 ;
        RECT 1758.965 4995.885 1836.970 4996.485 ;
        RECT 2303.965 4995.885 2381.970 4996.485 ;
        RECT 2848.965 4995.885 2922.035 4996.485 ;
        RECT 3388.000 4995.885 3435.335 4996.485 ;
        RECT 152.665 4992.185 202.330 4995.885 ;
        RECT 152.665 4990.000 186.065 4992.185 ;
        RECT 152.665 4989.875 169.115 4990.000 ;
        RECT 152.665 4988.000 153.365 4989.875 ;
        RECT 158.815 4989.785 169.115 4989.875 ;
        RECT 158.815 4989.735 164.265 4989.785 ;
        RECT 152.665 4457.330 153.365 4458.035 ;
      LAYER met4 ;
        RECT 153.765 4457.730 158.415 4989.475 ;
      LAYER met4 ;
        RECT 158.815 4988.000 159.415 4989.735 ;
        RECT 158.815 4457.330 159.415 4458.035 ;
      LAYER met4 ;
        RECT 159.815 4457.730 163.265 4989.335 ;
      LAYER met4 ;
        RECT 163.665 4988.000 164.265 4989.735 ;
        RECT 163.665 4457.330 164.265 4458.035 ;
      LAYER met4 ;
        RECT 164.665 4457.730 168.115 4989.385 ;
      LAYER met4 ;
        RECT 168.515 4988.000 169.115 4989.785 ;
        RECT 174.565 4989.925 186.065 4990.000 ;
        RECT 168.515 4457.330 169.115 4458.035 ;
      LAYER met4 ;
        RECT 169.515 4457.730 174.165 4989.600 ;
      LAYER met4 ;
        RECT 174.565 4988.000 175.165 4989.925 ;
        RECT 180.615 4989.870 186.065 4989.925 ;
        RECT 174.565 4457.330 175.165 4458.035 ;
      LAYER met4 ;
        RECT 175.565 4457.730 180.215 4989.525 ;
      LAYER met4 ;
        RECT 180.615 4988.000 181.215 4989.870 ;
      LAYER met4 ;
        RECT 181.615 4458.035 185.065 4989.470 ;
      LAYER met4 ;
        RECT 185.465 4988.000 186.065 4989.870 ;
        RECT 180.615 4457.635 181.215 4458.035 ;
        RECT 185.465 4457.635 186.065 4458.035 ;
      LAYER met4 ;
        RECT 186.465 4457.730 191.115 4991.785 ;
      LAYER met4 ;
        RECT 191.515 4990.750 202.330 4992.185 ;
        RECT 191.515 4988.000 192.115 4990.750 ;
        RECT 180.615 4457.330 186.065 4457.635 ;
        RECT 191.515 4457.330 192.115 4458.035 ;
      LAYER met4 ;
        RECT 192.515 4457.730 197.965 4990.350 ;
      LAYER met4 ;
        RECT 198.365 4989.635 202.330 4990.750 ;
      LAYER met4 ;
        RECT 202.730 4990.035 669.270 4995.485 ;
      LAYER met4 ;
        RECT 669.670 4989.635 746.330 4995.885 ;
      LAYER met4 ;
        RECT 746.730 4990.035 1214.270 4995.485 ;
      LAYER met4 ;
        RECT 1214.670 4989.635 1291.330 4995.885 ;
      LAYER met4 ;
        RECT 1291.730 4990.035 1759.270 4995.485 ;
      LAYER met4 ;
        RECT 1759.670 4989.635 1836.330 4995.885 ;
      LAYER met4 ;
        RECT 1836.730 4990.035 2304.270 4995.485 ;
      LAYER met4 ;
        RECT 2304.670 4989.635 2381.330 4995.885 ;
      LAYER met4 ;
        RECT 2381.730 4990.035 2849.270 4995.485 ;
      LAYER met4 ;
        RECT 2849.670 4990.035 2921.330 4995.885 ;
      LAYER met4 ;
        RECT 2921.730 4990.035 3390.350 4995.485 ;
      LAYER met4 ;
        RECT 3390.750 4989.635 3435.335 4995.885 ;
        RECT 198.365 4988.000 202.745 4989.635 ;
        RECT 668.965 4988.535 746.970 4989.635 ;
        RECT 1213.965 4988.535 1291.970 4989.635 ;
        RECT 1758.965 4988.535 1836.970 4989.635 ;
        RECT 2303.965 4988.535 2381.970 4989.635 ;
        RECT 3388.000 4985.670 3435.335 4989.635 ;
        RECT 3388.000 4985.255 3389.635 4985.670 ;
        RECT 152.665 4385.670 197.965 4457.330 ;
      LAYER met4 ;
        RECT 3390.035 4453.730 3395.485 4985.270 ;
      LAYER met4 ;
        RECT 3395.885 4985.255 3396.485 4985.670 ;
        RECT 3401.935 4985.655 3407.385 4985.670 ;
        RECT 3395.885 4453.330 3396.485 4454.035 ;
      LAYER met4 ;
        RECT 3396.885 4453.730 3401.535 4985.270 ;
      LAYER met4 ;
        RECT 3401.935 4985.255 3402.535 4985.655 ;
        RECT 3406.785 4985.255 3407.385 4985.655 ;
      LAYER met4 ;
        RECT 3402.935 4454.035 3406.385 4985.255 ;
      LAYER met4 ;
        RECT 3401.935 4453.635 3402.535 4454.035 ;
        RECT 3406.785 4453.635 3407.385 4454.035 ;
      LAYER met4 ;
        RECT 3407.785 4453.730 3412.435 4985.270 ;
      LAYER met4 ;
        RECT 3412.835 4985.255 3413.435 4985.670 ;
        RECT 3401.935 4453.330 3407.385 4453.635 ;
        RECT 3412.835 4453.330 3413.435 4454.035 ;
      LAYER met4 ;
        RECT 3413.835 4453.730 3418.485 4985.270 ;
      LAYER met4 ;
        RECT 3418.885 4985.255 3419.485 4985.670 ;
        RECT 3418.885 4453.330 3419.485 4454.035 ;
      LAYER met4 ;
        RECT 3419.885 4453.730 3423.335 4985.270 ;
      LAYER met4 ;
        RECT 3423.735 4985.255 3424.335 4985.670 ;
        RECT 3423.735 4453.330 3424.335 4454.035 ;
      LAYER met4 ;
        RECT 3424.735 4453.730 3428.185 4985.270 ;
      LAYER met4 ;
        RECT 3428.585 4985.255 3429.185 4985.670 ;
        RECT 3428.585 4453.330 3429.185 4454.035 ;
      LAYER met4 ;
        RECT 3429.585 4453.730 3434.235 4985.270 ;
      LAYER met4 ;
        RECT 3434.635 4985.255 3435.335 4985.670 ;
        RECT 3434.635 4453.330 3435.335 4454.035 ;
        RECT 152.665 4384.965 153.365 4385.670 ;
        RECT 152.665 3853.330 153.365 3853.970 ;
      LAYER met4 ;
        RECT 153.765 3853.730 158.415 4385.270 ;
      LAYER met4 ;
        RECT 158.815 4384.965 159.415 4385.670 ;
        RECT 158.815 3853.330 159.415 3853.970 ;
      LAYER met4 ;
        RECT 159.815 3853.730 163.265 4385.270 ;
      LAYER met4 ;
        RECT 163.665 4384.965 164.265 4385.670 ;
        RECT 163.665 3853.330 164.265 3853.970 ;
      LAYER met4 ;
        RECT 164.665 3853.730 168.115 4385.270 ;
      LAYER met4 ;
        RECT 168.515 4384.965 169.115 4385.670 ;
        RECT 168.515 3853.330 169.115 3853.970 ;
      LAYER met4 ;
        RECT 169.515 3853.730 174.165 4385.270 ;
      LAYER met4 ;
        RECT 174.565 4384.965 175.165 4385.670 ;
        RECT 180.615 4385.365 186.065 4385.670 ;
        RECT 174.565 3853.330 175.165 3853.970 ;
      LAYER met4 ;
        RECT 175.565 3853.730 180.215 4385.270 ;
      LAYER met4 ;
        RECT 180.615 4384.965 181.215 4385.365 ;
        RECT 185.465 4384.965 186.065 4385.365 ;
      LAYER met4 ;
        RECT 181.615 3853.970 185.065 4384.965 ;
      LAYER met4 ;
        RECT 180.615 3853.570 181.215 3853.970 ;
        RECT 185.465 3853.570 186.065 3853.970 ;
      LAYER met4 ;
        RECT 186.465 3853.730 191.115 4385.270 ;
      LAYER met4 ;
        RECT 191.515 4384.965 192.115 4385.670 ;
        RECT 180.615 3853.330 186.065 3853.570 ;
        RECT 191.515 3853.330 192.115 3853.970 ;
      LAYER met4 ;
        RECT 192.515 3853.730 197.965 4385.270 ;
      LAYER met4 ;
        RECT 3390.035 4381.670 3435.335 4453.330 ;
      LAYER met4 ;
        RECT 3387.735 4364.050 3388.065 4364.065 ;
        RECT 3382.230 4363.750 3388.065 4364.050 ;
        RECT 3382.230 4279.490 3382.530 4363.750 ;
        RECT 3387.735 4363.735 3388.065 4363.750 ;
        RECT 3381.790 4278.310 3382.970 4279.490 ;
        RECT 3380.870 4274.910 3382.050 4276.090 ;
        RECT 3381.310 4183.850 3381.610 4274.910 ;
        RECT 3381.310 4183.550 3382.530 4183.850 ;
        RECT 3382.230 4058.050 3382.530 4183.550 ;
        RECT 3382.230 4057.750 3383.450 4058.050 ;
        RECT 3383.150 3891.450 3383.450 4057.750 ;
        RECT 3381.310 3891.150 3383.450 3891.450 ;
      LAYER met4 ;
        RECT 198.365 3853.330 199.465 3853.970 ;
        RECT 152.665 3821.690 199.465 3853.330 ;
        RECT 152.035 3778.010 199.465 3821.690 ;
      LAYER met4 ;
        RECT 3381.310 3817.090 3381.610 3891.150 ;
      LAYER met4 ;
        RECT 3388.535 3849.330 3389.635 3850.035 ;
      LAYER met4 ;
        RECT 3390.035 3849.730 3395.485 4381.270 ;
      LAYER met4 ;
        RECT 3395.885 4380.965 3396.485 4381.670 ;
        RECT 3401.935 4381.365 3407.385 4381.670 ;
        RECT 3395.885 3849.330 3396.485 3850.035 ;
      LAYER met4 ;
        RECT 3396.885 3849.730 3401.535 4381.270 ;
      LAYER met4 ;
        RECT 3401.935 4380.965 3402.535 4381.365 ;
        RECT 3406.785 4380.965 3407.385 4381.365 ;
      LAYER met4 ;
        RECT 3402.935 3850.035 3406.385 4380.965 ;
      LAYER met4 ;
        RECT 3401.935 3849.635 3402.535 3850.035 ;
        RECT 3406.785 3849.635 3407.385 3850.035 ;
      LAYER met4 ;
        RECT 3407.785 3849.730 3412.435 4381.270 ;
      LAYER met4 ;
        RECT 3412.835 4380.965 3413.435 4381.670 ;
        RECT 3401.935 3849.330 3407.385 3849.635 ;
        RECT 3412.835 3849.330 3413.435 3850.035 ;
      LAYER met4 ;
        RECT 3413.835 3849.730 3418.485 4381.270 ;
      LAYER met4 ;
        RECT 3418.885 4380.965 3419.485 4381.670 ;
        RECT 3418.885 3849.330 3419.485 3850.035 ;
      LAYER met4 ;
        RECT 3419.885 3849.730 3423.335 4381.270 ;
      LAYER met4 ;
        RECT 3423.735 4380.965 3424.335 4381.670 ;
        RECT 3423.735 3849.330 3424.335 3850.035 ;
      LAYER met4 ;
        RECT 3424.735 3849.730 3428.185 4381.270 ;
      LAYER met4 ;
        RECT 3428.585 4380.965 3429.185 4381.670 ;
        RECT 3428.585 3849.330 3429.185 3850.035 ;
      LAYER met4 ;
        RECT 3429.585 3849.730 3434.235 4381.270 ;
      LAYER met4 ;
        RECT 3434.635 4380.965 3435.335 4381.670 ;
        RECT 3434.635 3849.330 3435.335 3850.035 ;
        RECT 3388.535 3847.990 3435.335 3849.330 ;
      LAYER met4 ;
        RECT 3435.735 3848.390 3436.065 5007.575 ;
      LAYER met4 ;
        RECT 3436.465 5005.955 3440.725 5007.975 ;
        RECT 3436.465 5005.275 3439.245 5005.955 ;
      LAYER met4 ;
        RECT 3380.870 3815.910 3382.050 3817.090 ;
        RECT 3386.390 3815.910 3387.570 3817.090 ;
      LAYER met4 ;
        RECT 147.275 3219.545 151.535 3221.065 ;
        RECT 147.275 3205.360 148.255 3219.545 ;
        RECT 0.000 3203.840 148.255 3205.360 ;
        RECT 0.000 3170.010 143.495 3203.840 ;
        RECT 0.000 3168.670 142.865 3170.010 ;
      LAYER met4 ;
        RECT 0.000 3167.000 24.215 3168.270 ;
      LAYER met4 ;
        RECT 24.615 3167.965 104.600 3168.670 ;
        RECT 0.000 2638.000 25.965 3167.000 ;
        RECT 102.965 3162.000 105.000 3167.000 ;
      LAYER met4 ;
        RECT 105.000 3162.000 129.965 3168.270 ;
      LAYER met4 ;
        RECT 130.365 3167.965 131.065 3168.670 ;
        RECT 129.965 3162.000 131.065 3167.000 ;
        RECT 102.965 3159.000 131.065 3162.000 ;
        RECT 102.965 3157.000 105.000 3159.000 ;
      LAYER met4 ;
        RECT 105.000 3157.000 129.965 3159.000 ;
      LAYER met4 ;
        RECT 129.965 3157.000 131.065 3159.000 ;
        RECT 102.965 3139.000 131.065 3157.000 ;
        RECT 102.965 3137.000 105.000 3139.000 ;
      LAYER met4 ;
        RECT 105.000 3137.000 129.965 3139.000 ;
      LAYER met4 ;
        RECT 129.965 3137.000 131.065 3139.000 ;
        RECT 102.965 3119.000 131.065 3137.000 ;
        RECT 102.965 3117.000 105.000 3119.000 ;
      LAYER met4 ;
        RECT 105.000 3117.000 129.965 3119.000 ;
      LAYER met4 ;
        RECT 129.965 3117.000 131.065 3119.000 ;
        RECT 102.965 3099.000 131.065 3117.000 ;
        RECT 102.965 3097.000 105.000 3099.000 ;
      LAYER met4 ;
        RECT 105.000 3097.000 129.965 3099.000 ;
      LAYER met4 ;
        RECT 129.965 3097.000 131.065 3099.000 ;
        RECT 102.965 3079.000 131.065 3097.000 ;
        RECT 102.965 3077.000 105.000 3079.000 ;
      LAYER met4 ;
        RECT 105.000 3077.000 129.965 3079.000 ;
      LAYER met4 ;
        RECT 129.965 3077.000 131.065 3079.000 ;
        RECT 102.965 3059.000 131.065 3077.000 ;
        RECT 102.965 3057.000 105.000 3059.000 ;
      LAYER met4 ;
        RECT 105.000 3057.000 129.965 3059.000 ;
      LAYER met4 ;
        RECT 129.965 3057.000 131.065 3059.000 ;
        RECT 102.965 3039.000 131.065 3057.000 ;
        RECT 102.965 3037.000 105.000 3039.000 ;
      LAYER met4 ;
        RECT 105.000 3037.000 129.965 3039.000 ;
      LAYER met4 ;
        RECT 129.965 3037.000 131.065 3039.000 ;
        RECT 102.965 3019.000 131.065 3037.000 ;
        RECT 102.965 3017.000 105.000 3019.000 ;
      LAYER met4 ;
        RECT 105.000 3017.000 129.965 3019.000 ;
      LAYER met4 ;
        RECT 129.965 3017.000 131.065 3019.000 ;
        RECT 102.965 2999.000 131.065 3017.000 ;
        RECT 102.965 2997.000 105.000 2999.000 ;
      LAYER met4 ;
        RECT 105.000 2997.000 129.965 2999.000 ;
      LAYER met4 ;
        RECT 129.965 2997.000 131.065 2999.000 ;
        RECT 102.965 2979.000 131.065 2997.000 ;
        RECT 102.965 2977.000 105.000 2979.000 ;
      LAYER met4 ;
        RECT 105.000 2977.000 129.965 2979.000 ;
      LAYER met4 ;
        RECT 129.965 2977.000 131.065 2979.000 ;
        RECT 102.965 2959.000 131.065 2977.000 ;
        RECT 102.965 2957.000 105.000 2959.000 ;
      LAYER met4 ;
        RECT 105.000 2957.000 129.965 2959.000 ;
      LAYER met4 ;
        RECT 129.965 2957.000 131.065 2959.000 ;
        RECT 102.965 2939.000 131.065 2957.000 ;
        RECT 102.965 2937.000 105.000 2939.000 ;
      LAYER met4 ;
        RECT 105.000 2937.000 129.965 2939.000 ;
      LAYER met4 ;
        RECT 129.965 2937.000 131.065 2939.000 ;
        RECT 102.965 2919.000 131.065 2937.000 ;
        RECT 102.965 2917.000 105.000 2919.000 ;
      LAYER met4 ;
        RECT 105.000 2917.000 129.965 2919.000 ;
      LAYER met4 ;
        RECT 129.965 2917.000 131.065 2919.000 ;
        RECT 102.965 2899.000 131.065 2917.000 ;
        RECT 102.965 2897.000 105.000 2899.000 ;
      LAYER met4 ;
        RECT 105.000 2897.000 129.965 2899.000 ;
      LAYER met4 ;
        RECT 129.965 2897.000 131.065 2899.000 ;
        RECT 102.965 2879.000 131.065 2897.000 ;
        RECT 102.965 2877.000 105.000 2879.000 ;
      LAYER met4 ;
        RECT 105.000 2877.000 129.965 2879.000 ;
      LAYER met4 ;
        RECT 129.965 2877.000 131.065 2879.000 ;
        RECT 102.965 2859.000 131.065 2877.000 ;
        RECT 102.965 2857.000 105.000 2859.000 ;
      LAYER met4 ;
        RECT 105.000 2857.000 129.965 2859.000 ;
      LAYER met4 ;
        RECT 129.965 2857.000 131.065 2859.000 ;
        RECT 102.965 2839.000 131.065 2857.000 ;
        RECT 102.965 2837.000 105.000 2839.000 ;
      LAYER met4 ;
        RECT 105.000 2837.000 129.965 2839.000 ;
      LAYER met4 ;
        RECT 129.965 2837.000 131.065 2839.000 ;
        RECT 102.965 2819.000 131.065 2837.000 ;
        RECT 102.965 2817.000 105.000 2819.000 ;
      LAYER met4 ;
        RECT 105.000 2817.000 129.965 2819.000 ;
      LAYER met4 ;
        RECT 129.965 2817.000 131.065 2819.000 ;
        RECT 102.965 2799.000 131.065 2817.000 ;
        RECT 102.965 2797.000 105.000 2799.000 ;
      LAYER met4 ;
        RECT 105.000 2797.000 129.965 2799.000 ;
      LAYER met4 ;
        RECT 129.965 2797.000 131.065 2799.000 ;
        RECT 102.965 2779.000 131.065 2797.000 ;
        RECT 102.965 2777.000 105.000 2779.000 ;
      LAYER met4 ;
        RECT 105.000 2777.000 129.965 2779.000 ;
      LAYER met4 ;
        RECT 129.965 2777.000 131.065 2779.000 ;
        RECT 102.965 2759.000 131.065 2777.000 ;
        RECT 102.965 2757.000 105.000 2759.000 ;
      LAYER met4 ;
        RECT 105.000 2757.000 129.965 2759.000 ;
      LAYER met4 ;
        RECT 129.965 2757.000 131.065 2759.000 ;
        RECT 102.965 2739.000 131.065 2757.000 ;
        RECT 102.965 2737.000 105.000 2739.000 ;
      LAYER met4 ;
        RECT 105.000 2737.000 129.965 2739.000 ;
      LAYER met4 ;
        RECT 129.965 2737.000 131.065 2739.000 ;
        RECT 102.965 2719.000 131.065 2737.000 ;
        RECT 102.965 2717.000 105.000 2719.000 ;
      LAYER met4 ;
        RECT 105.000 2717.000 129.965 2719.000 ;
      LAYER met4 ;
        RECT 129.965 2717.000 131.065 2719.000 ;
        RECT 102.965 2699.000 131.065 2717.000 ;
        RECT 102.965 2697.000 105.000 2699.000 ;
      LAYER met4 ;
        RECT 105.000 2697.000 129.965 2699.000 ;
      LAYER met4 ;
        RECT 129.965 2697.000 131.065 2699.000 ;
        RECT 102.965 2679.000 131.065 2697.000 ;
        RECT 102.965 2677.000 105.000 2679.000 ;
      LAYER met4 ;
        RECT 105.000 2677.000 129.965 2679.000 ;
      LAYER met4 ;
        RECT 129.965 2677.000 131.065 2679.000 ;
        RECT 102.965 2659.000 131.065 2677.000 ;
        RECT 102.965 2657.000 105.000 2659.000 ;
      LAYER met4 ;
        RECT 105.000 2657.000 129.965 2659.000 ;
      LAYER met4 ;
        RECT 129.965 2657.000 131.065 2659.000 ;
        RECT 102.965 2639.000 131.065 2657.000 ;
        RECT 102.965 2638.000 105.000 2639.000 ;
      LAYER met4 ;
        RECT 0.000 2636.730 24.215 2638.000 ;
      LAYER met4 ;
        RECT 24.615 2636.330 104.600 2636.970 ;
      LAYER met4 ;
        RECT 105.000 2636.730 129.965 2639.000 ;
      LAYER met4 ;
        RECT 129.965 2638.000 131.065 2639.000 ;
        RECT 130.365 2636.330 131.065 2636.970 ;
      LAYER met4 ;
        RECT 131.465 2636.730 135.915 3168.270 ;
      LAYER met4 ;
        RECT 136.315 3167.965 136.915 3168.670 ;
        RECT 136.315 2638.000 136.915 3163.000 ;
        RECT 136.315 2636.330 136.915 2636.970 ;
      LAYER met4 ;
        RECT 137.315 2636.730 141.765 3168.270 ;
      LAYER met4 ;
        RECT 142.165 3167.965 142.865 3168.670 ;
        RECT 142.165 2638.000 142.865 3167.000 ;
        RECT 142.165 2636.330 142.865 2636.970 ;
        RECT 0.000 2604.690 142.865 2636.330 ;
      LAYER met4 ;
        RECT 143.265 2605.090 143.595 3169.610 ;
      LAYER met4 ;
        RECT 0.000 2596.360 143.495 2604.690 ;
      LAYER met4 ;
        RECT 143.895 2596.760 146.875 3203.440 ;
      LAYER met4 ;
        RECT 147.275 3168.670 148.255 3203.840 ;
      LAYER met4 ;
        RECT 147.175 3167.000 148.355 3168.270 ;
      LAYER met4 ;
        RECT 147.275 2638.000 148.255 3167.000 ;
      LAYER met4 ;
        RECT 147.175 2636.730 148.355 2638.000 ;
      LAYER met4 ;
        RECT 147.275 2612.065 148.255 2636.330 ;
      LAYER met4 ;
        RECT 148.655 2612.465 151.635 3219.145 ;
        RECT 151.935 3214.090 152.265 3777.610 ;
      LAYER met4 ;
        RECT 152.665 3776.670 199.465 3778.010 ;
        RECT 152.665 3775.965 153.365 3776.670 ;
        RECT 152.665 3245.330 153.365 3245.970 ;
      LAYER met4 ;
        RECT 153.765 3245.730 158.415 3776.270 ;
      LAYER met4 ;
        RECT 158.815 3775.965 159.415 3776.670 ;
        RECT 158.815 3245.330 159.415 3245.970 ;
      LAYER met4 ;
        RECT 159.815 3245.730 163.265 3776.270 ;
      LAYER met4 ;
        RECT 163.665 3775.965 164.265 3776.670 ;
        RECT 163.665 3245.330 164.265 3245.970 ;
      LAYER met4 ;
        RECT 164.665 3245.730 168.115 3776.270 ;
      LAYER met4 ;
        RECT 168.515 3775.965 169.115 3776.670 ;
        RECT 168.515 3245.330 169.115 3245.970 ;
      LAYER met4 ;
        RECT 169.515 3245.730 174.165 3776.270 ;
      LAYER met4 ;
        RECT 174.565 3775.965 175.165 3776.670 ;
        RECT 180.615 3776.365 186.065 3776.670 ;
        RECT 174.565 3245.330 175.165 3245.970 ;
      LAYER met4 ;
        RECT 175.565 3245.730 180.215 3776.270 ;
      LAYER met4 ;
        RECT 180.615 3775.965 181.215 3776.365 ;
        RECT 185.465 3775.965 186.065 3776.365 ;
      LAYER met4 ;
        RECT 181.615 3245.970 185.065 3775.965 ;
      LAYER met4 ;
        RECT 180.615 3245.570 181.215 3245.970 ;
        RECT 185.465 3245.570 186.065 3245.970 ;
      LAYER met4 ;
        RECT 186.465 3245.730 191.115 3776.270 ;
      LAYER met4 ;
        RECT 191.515 3775.965 192.115 3776.670 ;
        RECT 180.615 3245.330 186.065 3245.570 ;
        RECT 191.515 3245.330 192.115 3245.970 ;
      LAYER met4 ;
        RECT 192.515 3245.730 197.965 3776.270 ;
      LAYER met4 ;
        RECT 198.365 3775.965 199.465 3776.670 ;
      LAYER met4 ;
        RECT 3386.830 3769.050 3387.130 3815.910 ;
      LAYER met4 ;
        RECT 3388.535 3804.310 3435.965 3847.990 ;
        RECT 3388.535 3772.670 3435.335 3804.310 ;
        RECT 3388.535 3772.030 3389.635 3772.670 ;
      LAYER met4 ;
        RECT 3383.150 3768.750 3387.130 3769.050 ;
        RECT 3383.150 3697.650 3383.450 3768.750 ;
        RECT 3383.150 3697.350 3384.370 3697.650 ;
        RECT 3384.070 3670.450 3384.370 3697.350 ;
        RECT 3384.070 3670.150 3386.210 3670.450 ;
        RECT 3385.910 3575.690 3386.210 3670.150 ;
        RECT 3382.710 3574.510 3383.890 3575.690 ;
        RECT 3385.470 3574.510 3386.650 3575.690 ;
        RECT 3383.150 3527.650 3383.450 3574.510 ;
        RECT 3383.150 3527.350 3384.370 3527.650 ;
        RECT 3384.070 3408.650 3384.370 3527.350 ;
        RECT 3383.150 3408.350 3384.370 3408.650 ;
        RECT 3383.150 3330.450 3383.450 3408.350 ;
        RECT 3382.230 3330.150 3383.450 3330.450 ;
      LAYER met4 ;
        RECT 198.365 3245.330 199.465 3245.970 ;
        RECT 152.665 3213.690 199.465 3245.330 ;
      LAYER met4 ;
        RECT 3382.230 3214.850 3382.530 3330.150 ;
      LAYER met4 ;
        RECT 3388.535 3241.330 3389.635 3242.035 ;
      LAYER met4 ;
        RECT 3390.035 3241.730 3395.485 3772.270 ;
      LAYER met4 ;
        RECT 3395.885 3772.030 3396.485 3772.670 ;
        RECT 3401.935 3772.430 3407.385 3772.670 ;
        RECT 3395.885 3241.330 3396.485 3242.035 ;
      LAYER met4 ;
        RECT 3396.885 3241.730 3401.535 3772.270 ;
      LAYER met4 ;
        RECT 3401.935 3772.030 3402.535 3772.430 ;
        RECT 3406.785 3772.030 3407.385 3772.430 ;
      LAYER met4 ;
        RECT 3402.935 3242.035 3406.385 3772.030 ;
      LAYER met4 ;
        RECT 3401.935 3241.635 3402.535 3242.035 ;
        RECT 3406.785 3241.635 3407.385 3242.035 ;
      LAYER met4 ;
        RECT 3407.785 3241.730 3412.435 3772.270 ;
      LAYER met4 ;
        RECT 3412.835 3772.030 3413.435 3772.670 ;
        RECT 3401.935 3241.330 3407.385 3241.635 ;
        RECT 3412.835 3241.330 3413.435 3242.035 ;
      LAYER met4 ;
        RECT 3413.835 3241.730 3418.485 3772.270 ;
      LAYER met4 ;
        RECT 3418.885 3772.030 3419.485 3772.670 ;
        RECT 3418.885 3241.330 3419.485 3242.035 ;
      LAYER met4 ;
        RECT 3419.885 3241.730 3423.335 3772.270 ;
      LAYER met4 ;
        RECT 3423.735 3772.030 3424.335 3772.670 ;
        RECT 3423.735 3241.330 3424.335 3242.035 ;
      LAYER met4 ;
        RECT 3424.735 3241.730 3428.185 3772.270 ;
      LAYER met4 ;
        RECT 3428.585 3772.030 3429.185 3772.670 ;
        RECT 3428.585 3241.330 3429.185 3242.035 ;
      LAYER met4 ;
        RECT 3429.585 3241.730 3434.235 3772.270 ;
      LAYER met4 ;
        RECT 3434.635 3772.030 3435.335 3772.670 ;
        RECT 3434.635 3241.330 3435.335 3242.035 ;
        RECT 3388.535 3239.990 3435.335 3241.330 ;
      LAYER met4 ;
        RECT 3435.735 3240.390 3436.065 3803.910 ;
        RECT 3436.365 3798.855 3439.345 5004.875 ;
        RECT 3439.645 4984.000 3440.825 5005.555 ;
      LAYER met4 ;
        RECT 3439.745 4455.000 3440.725 4984.000 ;
      LAYER met4 ;
        RECT 3439.645 4453.730 3440.825 4455.000 ;
      LAYER met4 ;
        RECT 3439.745 4381.670 3440.725 4453.330 ;
      LAYER met4 ;
        RECT 3439.645 4380.000 3440.825 4381.270 ;
      LAYER met4 ;
        RECT 3439.745 3851.000 3440.725 4380.000 ;
      LAYER met4 ;
        RECT 3439.645 3849.730 3440.825 3851.000 ;
      LAYER met4 ;
        RECT 3439.745 3814.160 3440.725 3849.330 ;
      LAYER met4 ;
        RECT 3441.125 3814.560 3444.105 5010.910 ;
        RECT 3444.405 3848.390 3444.735 5011.175 ;
      LAYER met4 ;
        RECT 3445.135 4986.255 3588.000 5011.575 ;
        RECT 3445.135 4985.670 3457.635 4986.255 ;
        RECT 3445.135 4985.255 3445.835 4985.670 ;
        RECT 3445.135 4455.000 3445.835 4984.000 ;
        RECT 3445.135 4453.330 3445.835 4454.035 ;
      LAYER met4 ;
        RECT 3446.235 4453.730 3450.685 4985.270 ;
      LAYER met4 ;
        RECT 3451.085 4985.255 3451.685 4985.670 ;
        RECT 3451.085 4455.000 3451.685 4980.000 ;
        RECT 3451.085 4453.330 3451.685 4454.035 ;
      LAYER met4 ;
        RECT 3452.085 4453.730 3456.535 4985.270 ;
      LAYER met4 ;
        RECT 3456.935 4985.255 3457.635 4985.670 ;
        RECT 3456.935 4979.000 3458.035 4984.000 ;
      LAYER met4 ;
        RECT 3458.035 4979.000 3483.000 4985.855 ;
      LAYER met4 ;
        RECT 3483.400 4985.670 3588.000 4986.255 ;
        RECT 3483.400 4985.255 3563.385 4985.670 ;
      LAYER met4 ;
        RECT 3563.785 4984.000 3588.000 4985.270 ;
      LAYER met4 ;
        RECT 3483.000 4979.000 3485.035 4984.000 ;
        RECT 3456.935 4976.000 3485.035 4979.000 ;
        RECT 3456.935 4974.000 3458.035 4976.000 ;
      LAYER met4 ;
        RECT 3458.035 4974.000 3483.000 4976.000 ;
      LAYER met4 ;
        RECT 3483.000 4974.000 3485.035 4976.000 ;
        RECT 3456.935 4956.000 3485.035 4974.000 ;
        RECT 3456.935 4954.000 3458.035 4956.000 ;
      LAYER met4 ;
        RECT 3458.035 4954.000 3483.000 4956.000 ;
      LAYER met4 ;
        RECT 3483.000 4954.000 3485.035 4956.000 ;
        RECT 3456.935 4936.000 3485.035 4954.000 ;
        RECT 3456.935 4934.000 3458.035 4936.000 ;
      LAYER met4 ;
        RECT 3458.035 4934.000 3483.000 4936.000 ;
      LAYER met4 ;
        RECT 3483.000 4934.000 3485.035 4936.000 ;
        RECT 3456.935 4916.000 3485.035 4934.000 ;
        RECT 3456.935 4914.000 3458.035 4916.000 ;
      LAYER met4 ;
        RECT 3458.035 4914.000 3483.000 4916.000 ;
      LAYER met4 ;
        RECT 3483.000 4914.000 3485.035 4916.000 ;
        RECT 3456.935 4896.000 3485.035 4914.000 ;
        RECT 3456.935 4894.000 3458.035 4896.000 ;
      LAYER met4 ;
        RECT 3458.035 4894.000 3483.000 4896.000 ;
      LAYER met4 ;
        RECT 3483.000 4894.000 3485.035 4896.000 ;
        RECT 3456.935 4876.000 3485.035 4894.000 ;
        RECT 3456.935 4874.000 3458.035 4876.000 ;
      LAYER met4 ;
        RECT 3458.035 4874.000 3483.000 4876.000 ;
      LAYER met4 ;
        RECT 3483.000 4874.000 3485.035 4876.000 ;
        RECT 3456.935 4856.000 3485.035 4874.000 ;
        RECT 3456.935 4854.000 3458.035 4856.000 ;
      LAYER met4 ;
        RECT 3458.035 4854.000 3483.000 4856.000 ;
      LAYER met4 ;
        RECT 3483.000 4854.000 3485.035 4856.000 ;
        RECT 3456.935 4836.000 3485.035 4854.000 ;
        RECT 3456.935 4834.000 3458.035 4836.000 ;
      LAYER met4 ;
        RECT 3458.035 4834.000 3483.000 4836.000 ;
      LAYER met4 ;
        RECT 3483.000 4834.000 3485.035 4836.000 ;
        RECT 3456.935 4816.000 3485.035 4834.000 ;
        RECT 3456.935 4814.000 3458.035 4816.000 ;
      LAYER met4 ;
        RECT 3458.035 4814.000 3483.000 4816.000 ;
      LAYER met4 ;
        RECT 3483.000 4814.000 3485.035 4816.000 ;
        RECT 3456.935 4796.000 3485.035 4814.000 ;
        RECT 3456.935 4794.000 3458.035 4796.000 ;
      LAYER met4 ;
        RECT 3458.035 4794.000 3483.000 4796.000 ;
      LAYER met4 ;
        RECT 3483.000 4794.000 3485.035 4796.000 ;
        RECT 3456.935 4776.000 3485.035 4794.000 ;
        RECT 3456.935 4774.000 3458.035 4776.000 ;
      LAYER met4 ;
        RECT 3458.035 4774.000 3483.000 4776.000 ;
      LAYER met4 ;
        RECT 3483.000 4774.000 3485.035 4776.000 ;
        RECT 3456.935 4756.000 3485.035 4774.000 ;
        RECT 3456.935 4754.000 3458.035 4756.000 ;
      LAYER met4 ;
        RECT 3458.035 4754.000 3483.000 4756.000 ;
      LAYER met4 ;
        RECT 3483.000 4754.000 3485.035 4756.000 ;
        RECT 3456.935 4736.000 3485.035 4754.000 ;
        RECT 3456.935 4734.000 3458.035 4736.000 ;
      LAYER met4 ;
        RECT 3458.035 4734.000 3483.000 4736.000 ;
      LAYER met4 ;
        RECT 3483.000 4734.000 3485.035 4736.000 ;
        RECT 3456.935 4716.000 3485.035 4734.000 ;
        RECT 3456.935 4714.000 3458.035 4716.000 ;
      LAYER met4 ;
        RECT 3458.035 4714.000 3483.000 4716.000 ;
      LAYER met4 ;
        RECT 3483.000 4714.000 3485.035 4716.000 ;
        RECT 3456.935 4696.000 3485.035 4714.000 ;
        RECT 3456.935 4694.000 3458.035 4696.000 ;
      LAYER met4 ;
        RECT 3458.035 4694.000 3483.000 4696.000 ;
      LAYER met4 ;
        RECT 3483.000 4694.000 3485.035 4696.000 ;
        RECT 3456.935 4676.000 3485.035 4694.000 ;
        RECT 3456.935 4674.000 3458.035 4676.000 ;
      LAYER met4 ;
        RECT 3458.035 4674.000 3483.000 4676.000 ;
      LAYER met4 ;
        RECT 3483.000 4674.000 3485.035 4676.000 ;
        RECT 3456.935 4656.000 3485.035 4674.000 ;
        RECT 3456.935 4654.000 3458.035 4656.000 ;
      LAYER met4 ;
        RECT 3458.035 4654.000 3483.000 4656.000 ;
      LAYER met4 ;
        RECT 3483.000 4654.000 3485.035 4656.000 ;
        RECT 3456.935 4636.000 3485.035 4654.000 ;
        RECT 3456.935 4634.000 3458.035 4636.000 ;
      LAYER met4 ;
        RECT 3458.035 4634.000 3483.000 4636.000 ;
      LAYER met4 ;
        RECT 3483.000 4634.000 3485.035 4636.000 ;
        RECT 3456.935 4616.000 3485.035 4634.000 ;
        RECT 3456.935 4614.000 3458.035 4616.000 ;
      LAYER met4 ;
        RECT 3458.035 4614.000 3483.000 4616.000 ;
      LAYER met4 ;
        RECT 3483.000 4614.000 3485.035 4616.000 ;
        RECT 3456.935 4596.000 3485.035 4614.000 ;
        RECT 3456.935 4594.000 3458.035 4596.000 ;
      LAYER met4 ;
        RECT 3458.035 4594.000 3483.000 4596.000 ;
      LAYER met4 ;
        RECT 3483.000 4594.000 3485.035 4596.000 ;
        RECT 3456.935 4576.000 3485.035 4594.000 ;
        RECT 3456.935 4574.000 3458.035 4576.000 ;
      LAYER met4 ;
        RECT 3458.035 4574.000 3483.000 4576.000 ;
      LAYER met4 ;
        RECT 3483.000 4574.000 3485.035 4576.000 ;
        RECT 3456.935 4556.000 3485.035 4574.000 ;
        RECT 3456.935 4554.000 3458.035 4556.000 ;
      LAYER met4 ;
        RECT 3458.035 4554.000 3483.000 4556.000 ;
      LAYER met4 ;
        RECT 3483.000 4554.000 3485.035 4556.000 ;
        RECT 3456.935 4536.000 3485.035 4554.000 ;
        RECT 3456.935 4534.000 3458.035 4536.000 ;
      LAYER met4 ;
        RECT 3458.035 4534.000 3483.000 4536.000 ;
      LAYER met4 ;
        RECT 3483.000 4534.000 3485.035 4536.000 ;
        RECT 3456.935 4516.000 3485.035 4534.000 ;
        RECT 3456.935 4514.000 3458.035 4516.000 ;
      LAYER met4 ;
        RECT 3458.035 4514.000 3483.000 4516.000 ;
      LAYER met4 ;
        RECT 3483.000 4514.000 3485.035 4516.000 ;
        RECT 3456.935 4496.000 3485.035 4514.000 ;
        RECT 3456.935 4494.000 3458.035 4496.000 ;
      LAYER met4 ;
        RECT 3458.035 4494.000 3483.000 4496.000 ;
      LAYER met4 ;
        RECT 3483.000 4494.000 3485.035 4496.000 ;
        RECT 3456.935 4476.000 3485.035 4494.000 ;
        RECT 3456.935 4474.000 3458.035 4476.000 ;
      LAYER met4 ;
        RECT 3458.035 4474.000 3483.000 4476.000 ;
      LAYER met4 ;
        RECT 3483.000 4474.000 3485.035 4476.000 ;
        RECT 3456.935 4456.000 3485.035 4474.000 ;
        RECT 3456.935 4455.000 3458.035 4456.000 ;
        RECT 3456.935 4453.330 3457.635 4454.035 ;
      LAYER met4 ;
        RECT 3458.035 4453.730 3483.000 4456.000 ;
      LAYER met4 ;
        RECT 3483.000 4455.000 3485.035 4456.000 ;
        RECT 3562.035 4455.000 3588.000 4984.000 ;
        RECT 3483.400 4453.330 3563.385 4454.035 ;
      LAYER met4 ;
        RECT 3563.785 4453.730 3588.000 4455.000 ;
      LAYER met4 ;
        RECT 3445.135 4381.670 3588.000 4453.330 ;
        RECT 3445.135 4380.965 3445.835 4381.670 ;
        RECT 3445.135 3851.000 3445.835 4380.000 ;
        RECT 3445.135 3849.330 3445.835 3850.035 ;
      LAYER met4 ;
        RECT 3446.235 3849.730 3450.685 4381.270 ;
      LAYER met4 ;
        RECT 3451.085 4380.965 3451.685 4381.670 ;
        RECT 3451.085 3851.000 3451.685 4376.000 ;
        RECT 3451.085 3849.330 3451.685 3850.035 ;
      LAYER met4 ;
        RECT 3452.085 3849.730 3456.535 4381.270 ;
      LAYER met4 ;
        RECT 3456.935 4380.965 3457.635 4381.670 ;
        RECT 3456.935 4375.000 3458.035 4380.000 ;
      LAYER met4 ;
        RECT 3458.035 4375.000 3483.000 4381.270 ;
      LAYER met4 ;
        RECT 3483.400 4380.965 3563.385 4381.670 ;
      LAYER met4 ;
        RECT 3563.785 4380.000 3588.000 4381.270 ;
      LAYER met4 ;
        RECT 3483.000 4375.000 3485.035 4380.000 ;
        RECT 3456.935 4372.000 3485.035 4375.000 ;
        RECT 3456.935 4370.000 3458.035 4372.000 ;
      LAYER met4 ;
        RECT 3458.035 4370.000 3483.000 4372.000 ;
      LAYER met4 ;
        RECT 3483.000 4370.000 3485.035 4372.000 ;
        RECT 3456.935 4352.000 3485.035 4370.000 ;
        RECT 3456.935 4350.000 3458.035 4352.000 ;
      LAYER met4 ;
        RECT 3458.035 4350.000 3483.000 4352.000 ;
      LAYER met4 ;
        RECT 3483.000 4350.000 3485.035 4352.000 ;
        RECT 3456.935 4332.000 3485.035 4350.000 ;
        RECT 3456.935 4330.000 3458.035 4332.000 ;
      LAYER met4 ;
        RECT 3458.035 4330.000 3483.000 4332.000 ;
      LAYER met4 ;
        RECT 3483.000 4330.000 3485.035 4332.000 ;
        RECT 3456.935 4312.000 3485.035 4330.000 ;
        RECT 3456.935 4310.000 3458.035 4312.000 ;
      LAYER met4 ;
        RECT 3458.035 4310.000 3483.000 4312.000 ;
      LAYER met4 ;
        RECT 3483.000 4310.000 3485.035 4312.000 ;
        RECT 3456.935 4292.000 3485.035 4310.000 ;
        RECT 3456.935 4290.000 3458.035 4292.000 ;
      LAYER met4 ;
        RECT 3458.035 4290.000 3483.000 4292.000 ;
      LAYER met4 ;
        RECT 3483.000 4290.000 3485.035 4292.000 ;
        RECT 3456.935 4272.000 3485.035 4290.000 ;
        RECT 3456.935 4270.000 3458.035 4272.000 ;
      LAYER met4 ;
        RECT 3458.035 4270.000 3483.000 4272.000 ;
      LAYER met4 ;
        RECT 3483.000 4270.000 3485.035 4272.000 ;
        RECT 3456.935 4252.000 3485.035 4270.000 ;
        RECT 3456.935 4250.000 3458.035 4252.000 ;
      LAYER met4 ;
        RECT 3458.035 4250.000 3483.000 4252.000 ;
      LAYER met4 ;
        RECT 3483.000 4250.000 3485.035 4252.000 ;
        RECT 3456.935 4232.000 3485.035 4250.000 ;
        RECT 3456.935 4230.000 3458.035 4232.000 ;
      LAYER met4 ;
        RECT 3458.035 4230.000 3483.000 4232.000 ;
      LAYER met4 ;
        RECT 3483.000 4230.000 3485.035 4232.000 ;
        RECT 3456.935 4212.000 3485.035 4230.000 ;
        RECT 3456.935 4210.000 3458.035 4212.000 ;
      LAYER met4 ;
        RECT 3458.035 4210.000 3483.000 4212.000 ;
      LAYER met4 ;
        RECT 3483.000 4210.000 3485.035 4212.000 ;
        RECT 3456.935 4192.000 3485.035 4210.000 ;
        RECT 3456.935 4190.000 3458.035 4192.000 ;
      LAYER met4 ;
        RECT 3458.035 4190.000 3483.000 4192.000 ;
      LAYER met4 ;
        RECT 3483.000 4190.000 3485.035 4192.000 ;
        RECT 3456.935 4172.000 3485.035 4190.000 ;
        RECT 3456.935 4170.000 3458.035 4172.000 ;
      LAYER met4 ;
        RECT 3458.035 4170.000 3483.000 4172.000 ;
      LAYER met4 ;
        RECT 3483.000 4170.000 3485.035 4172.000 ;
        RECT 3456.935 4152.000 3485.035 4170.000 ;
        RECT 3456.935 4150.000 3458.035 4152.000 ;
      LAYER met4 ;
        RECT 3458.035 4150.000 3483.000 4152.000 ;
      LAYER met4 ;
        RECT 3483.000 4150.000 3485.035 4152.000 ;
        RECT 3456.935 4132.000 3485.035 4150.000 ;
        RECT 3456.935 4130.000 3458.035 4132.000 ;
      LAYER met4 ;
        RECT 3458.035 4130.000 3483.000 4132.000 ;
      LAYER met4 ;
        RECT 3483.000 4130.000 3485.035 4132.000 ;
        RECT 3456.935 4112.000 3485.035 4130.000 ;
        RECT 3456.935 4110.000 3458.035 4112.000 ;
      LAYER met4 ;
        RECT 3458.035 4110.000 3483.000 4112.000 ;
      LAYER met4 ;
        RECT 3483.000 4110.000 3485.035 4112.000 ;
        RECT 3456.935 4092.000 3485.035 4110.000 ;
        RECT 3456.935 4090.000 3458.035 4092.000 ;
      LAYER met4 ;
        RECT 3458.035 4090.000 3483.000 4092.000 ;
      LAYER met4 ;
        RECT 3483.000 4090.000 3485.035 4092.000 ;
        RECT 3456.935 4072.000 3485.035 4090.000 ;
        RECT 3456.935 4070.000 3458.035 4072.000 ;
      LAYER met4 ;
        RECT 3458.035 4070.000 3483.000 4072.000 ;
      LAYER met4 ;
        RECT 3483.000 4070.000 3485.035 4072.000 ;
        RECT 3456.935 4052.000 3485.035 4070.000 ;
        RECT 3456.935 4050.000 3458.035 4052.000 ;
      LAYER met4 ;
        RECT 3458.035 4050.000 3483.000 4052.000 ;
      LAYER met4 ;
        RECT 3483.000 4050.000 3485.035 4052.000 ;
        RECT 3456.935 4032.000 3485.035 4050.000 ;
        RECT 3456.935 4030.000 3458.035 4032.000 ;
      LAYER met4 ;
        RECT 3458.035 4030.000 3483.000 4032.000 ;
      LAYER met4 ;
        RECT 3483.000 4030.000 3485.035 4032.000 ;
        RECT 3456.935 4012.000 3485.035 4030.000 ;
        RECT 3456.935 4010.000 3458.035 4012.000 ;
      LAYER met4 ;
        RECT 3458.035 4010.000 3483.000 4012.000 ;
      LAYER met4 ;
        RECT 3483.000 4010.000 3485.035 4012.000 ;
        RECT 3456.935 3992.000 3485.035 4010.000 ;
        RECT 3456.935 3990.000 3458.035 3992.000 ;
      LAYER met4 ;
        RECT 3458.035 3990.000 3483.000 3992.000 ;
      LAYER met4 ;
        RECT 3483.000 3990.000 3485.035 3992.000 ;
        RECT 3456.935 3972.000 3485.035 3990.000 ;
        RECT 3456.935 3970.000 3458.035 3972.000 ;
      LAYER met4 ;
        RECT 3458.035 3970.000 3483.000 3972.000 ;
      LAYER met4 ;
        RECT 3483.000 3970.000 3485.035 3972.000 ;
        RECT 3456.935 3952.000 3485.035 3970.000 ;
        RECT 3456.935 3950.000 3458.035 3952.000 ;
      LAYER met4 ;
        RECT 3458.035 3950.000 3483.000 3952.000 ;
      LAYER met4 ;
        RECT 3483.000 3950.000 3485.035 3952.000 ;
        RECT 3456.935 3932.000 3485.035 3950.000 ;
        RECT 3456.935 3930.000 3458.035 3932.000 ;
      LAYER met4 ;
        RECT 3458.035 3930.000 3483.000 3932.000 ;
      LAYER met4 ;
        RECT 3483.000 3930.000 3485.035 3932.000 ;
        RECT 3456.935 3912.000 3485.035 3930.000 ;
        RECT 3456.935 3910.000 3458.035 3912.000 ;
      LAYER met4 ;
        RECT 3458.035 3910.000 3483.000 3912.000 ;
      LAYER met4 ;
        RECT 3483.000 3910.000 3485.035 3912.000 ;
        RECT 3456.935 3892.000 3485.035 3910.000 ;
        RECT 3456.935 3890.000 3458.035 3892.000 ;
      LAYER met4 ;
        RECT 3458.035 3890.000 3483.000 3892.000 ;
      LAYER met4 ;
        RECT 3483.000 3890.000 3485.035 3892.000 ;
        RECT 3456.935 3872.000 3485.035 3890.000 ;
        RECT 3456.935 3870.000 3458.035 3872.000 ;
      LAYER met4 ;
        RECT 3458.035 3870.000 3483.000 3872.000 ;
      LAYER met4 ;
        RECT 3483.000 3870.000 3485.035 3872.000 ;
        RECT 3456.935 3852.000 3485.035 3870.000 ;
        RECT 3456.935 3851.000 3458.035 3852.000 ;
        RECT 3456.935 3849.330 3457.635 3850.035 ;
      LAYER met4 ;
        RECT 3458.035 3849.730 3483.000 3852.000 ;
      LAYER met4 ;
        RECT 3483.000 3851.000 3485.035 3852.000 ;
        RECT 3562.035 3851.000 3588.000 4380.000 ;
        RECT 3483.400 3849.330 3563.385 3850.035 ;
      LAYER met4 ;
        RECT 3563.785 3849.730 3588.000 3851.000 ;
      LAYER met4 ;
        RECT 3445.135 3847.990 3588.000 3849.330 ;
        RECT 3444.505 3814.160 3588.000 3847.990 ;
        RECT 3439.745 3812.640 3588.000 3814.160 ;
        RECT 3439.745 3798.455 3440.725 3812.640 ;
        RECT 3436.465 3796.935 3440.725 3798.455 ;
      LAYER met4 ;
        RECT 3382.230 3214.550 3383.450 3214.850 ;
      LAYER met4 ;
        RECT 152.035 3170.010 199.465 3213.690 ;
        RECT 147.275 2610.545 151.535 2612.065 ;
        RECT 147.275 2596.360 148.255 2610.545 ;
        RECT 0.000 2594.840 148.255 2596.360 ;
        RECT 0.000 2561.010 143.495 2594.840 ;
        RECT 0.000 2559.670 142.865 2561.010 ;
      LAYER met4 ;
        RECT 0.000 2558.000 24.215 2559.270 ;
      LAYER met4 ;
        RECT 24.615 2558.965 104.600 2559.670 ;
        RECT 0.000 2029.000 25.965 2558.000 ;
        RECT 102.965 2553.000 105.000 2558.000 ;
      LAYER met4 ;
        RECT 105.000 2553.000 129.965 2559.270 ;
      LAYER met4 ;
        RECT 130.365 2558.965 131.065 2559.670 ;
        RECT 129.965 2553.000 131.065 2558.000 ;
        RECT 102.965 2550.000 131.065 2553.000 ;
        RECT 102.965 2548.000 105.000 2550.000 ;
      LAYER met4 ;
        RECT 105.000 2548.000 129.965 2550.000 ;
      LAYER met4 ;
        RECT 129.965 2548.000 131.065 2550.000 ;
        RECT 102.965 2530.000 131.065 2548.000 ;
        RECT 102.965 2528.000 105.000 2530.000 ;
      LAYER met4 ;
        RECT 105.000 2528.000 129.965 2530.000 ;
      LAYER met4 ;
        RECT 129.965 2528.000 131.065 2530.000 ;
        RECT 102.965 2510.000 131.065 2528.000 ;
        RECT 102.965 2508.000 105.000 2510.000 ;
      LAYER met4 ;
        RECT 105.000 2508.000 129.965 2510.000 ;
      LAYER met4 ;
        RECT 129.965 2508.000 131.065 2510.000 ;
        RECT 102.965 2490.000 131.065 2508.000 ;
        RECT 102.965 2488.000 105.000 2490.000 ;
      LAYER met4 ;
        RECT 105.000 2488.000 129.965 2490.000 ;
      LAYER met4 ;
        RECT 129.965 2488.000 131.065 2490.000 ;
        RECT 102.965 2470.000 131.065 2488.000 ;
        RECT 102.965 2468.000 105.000 2470.000 ;
      LAYER met4 ;
        RECT 105.000 2468.000 129.965 2470.000 ;
      LAYER met4 ;
        RECT 129.965 2468.000 131.065 2470.000 ;
        RECT 102.965 2450.000 131.065 2468.000 ;
        RECT 102.965 2448.000 105.000 2450.000 ;
      LAYER met4 ;
        RECT 105.000 2448.000 129.965 2450.000 ;
      LAYER met4 ;
        RECT 129.965 2448.000 131.065 2450.000 ;
        RECT 102.965 2430.000 131.065 2448.000 ;
        RECT 102.965 2428.000 105.000 2430.000 ;
      LAYER met4 ;
        RECT 105.000 2428.000 129.965 2430.000 ;
      LAYER met4 ;
        RECT 129.965 2428.000 131.065 2430.000 ;
        RECT 102.965 2410.000 131.065 2428.000 ;
        RECT 102.965 2408.000 105.000 2410.000 ;
      LAYER met4 ;
        RECT 105.000 2408.000 129.965 2410.000 ;
      LAYER met4 ;
        RECT 129.965 2408.000 131.065 2410.000 ;
        RECT 102.965 2390.000 131.065 2408.000 ;
        RECT 102.965 2388.000 105.000 2390.000 ;
      LAYER met4 ;
        RECT 105.000 2388.000 129.965 2390.000 ;
      LAYER met4 ;
        RECT 129.965 2388.000 131.065 2390.000 ;
        RECT 102.965 2370.000 131.065 2388.000 ;
        RECT 102.965 2368.000 105.000 2370.000 ;
      LAYER met4 ;
        RECT 105.000 2368.000 129.965 2370.000 ;
      LAYER met4 ;
        RECT 129.965 2368.000 131.065 2370.000 ;
        RECT 102.965 2350.000 131.065 2368.000 ;
        RECT 102.965 2348.000 105.000 2350.000 ;
      LAYER met4 ;
        RECT 105.000 2348.000 129.965 2350.000 ;
      LAYER met4 ;
        RECT 129.965 2348.000 131.065 2350.000 ;
        RECT 102.965 2330.000 131.065 2348.000 ;
        RECT 102.965 2328.000 105.000 2330.000 ;
      LAYER met4 ;
        RECT 105.000 2328.000 129.965 2330.000 ;
      LAYER met4 ;
        RECT 129.965 2328.000 131.065 2330.000 ;
        RECT 102.965 2310.000 131.065 2328.000 ;
        RECT 102.965 2308.000 105.000 2310.000 ;
      LAYER met4 ;
        RECT 105.000 2308.000 129.965 2310.000 ;
      LAYER met4 ;
        RECT 129.965 2308.000 131.065 2310.000 ;
        RECT 102.965 2290.000 131.065 2308.000 ;
        RECT 102.965 2288.000 105.000 2290.000 ;
      LAYER met4 ;
        RECT 105.000 2288.000 129.965 2290.000 ;
      LAYER met4 ;
        RECT 129.965 2288.000 131.065 2290.000 ;
        RECT 102.965 2270.000 131.065 2288.000 ;
        RECT 102.965 2268.000 105.000 2270.000 ;
      LAYER met4 ;
        RECT 105.000 2268.000 129.965 2270.000 ;
      LAYER met4 ;
        RECT 129.965 2268.000 131.065 2270.000 ;
        RECT 102.965 2250.000 131.065 2268.000 ;
        RECT 102.965 2248.000 105.000 2250.000 ;
      LAYER met4 ;
        RECT 105.000 2248.000 129.965 2250.000 ;
      LAYER met4 ;
        RECT 129.965 2248.000 131.065 2250.000 ;
        RECT 102.965 2230.000 131.065 2248.000 ;
        RECT 102.965 2228.000 105.000 2230.000 ;
      LAYER met4 ;
        RECT 105.000 2228.000 129.965 2230.000 ;
      LAYER met4 ;
        RECT 129.965 2228.000 131.065 2230.000 ;
        RECT 102.965 2210.000 131.065 2228.000 ;
        RECT 102.965 2208.000 105.000 2210.000 ;
      LAYER met4 ;
        RECT 105.000 2208.000 129.965 2210.000 ;
      LAYER met4 ;
        RECT 129.965 2208.000 131.065 2210.000 ;
        RECT 102.965 2190.000 131.065 2208.000 ;
        RECT 102.965 2188.000 105.000 2190.000 ;
      LAYER met4 ;
        RECT 105.000 2188.000 129.965 2190.000 ;
      LAYER met4 ;
        RECT 129.965 2188.000 131.065 2190.000 ;
        RECT 102.965 2170.000 131.065 2188.000 ;
        RECT 102.965 2168.000 105.000 2170.000 ;
      LAYER met4 ;
        RECT 105.000 2168.000 129.965 2170.000 ;
      LAYER met4 ;
        RECT 129.965 2168.000 131.065 2170.000 ;
        RECT 102.965 2150.000 131.065 2168.000 ;
        RECT 102.965 2148.000 105.000 2150.000 ;
      LAYER met4 ;
        RECT 105.000 2148.000 129.965 2150.000 ;
      LAYER met4 ;
        RECT 129.965 2148.000 131.065 2150.000 ;
        RECT 102.965 2130.000 131.065 2148.000 ;
        RECT 102.965 2128.000 105.000 2130.000 ;
      LAYER met4 ;
        RECT 105.000 2128.000 129.965 2130.000 ;
      LAYER met4 ;
        RECT 129.965 2128.000 131.065 2130.000 ;
        RECT 102.965 2110.000 131.065 2128.000 ;
        RECT 102.965 2108.000 105.000 2110.000 ;
      LAYER met4 ;
        RECT 105.000 2108.000 129.965 2110.000 ;
      LAYER met4 ;
        RECT 129.965 2108.000 131.065 2110.000 ;
        RECT 102.965 2090.000 131.065 2108.000 ;
        RECT 102.965 2088.000 105.000 2090.000 ;
      LAYER met4 ;
        RECT 105.000 2088.000 129.965 2090.000 ;
      LAYER met4 ;
        RECT 129.965 2088.000 131.065 2090.000 ;
        RECT 102.965 2070.000 131.065 2088.000 ;
        RECT 102.965 2068.000 105.000 2070.000 ;
      LAYER met4 ;
        RECT 105.000 2068.000 129.965 2070.000 ;
      LAYER met4 ;
        RECT 129.965 2068.000 131.065 2070.000 ;
        RECT 102.965 2050.000 131.065 2068.000 ;
        RECT 102.965 2048.000 105.000 2050.000 ;
      LAYER met4 ;
        RECT 105.000 2048.000 129.965 2050.000 ;
      LAYER met4 ;
        RECT 129.965 2048.000 131.065 2050.000 ;
        RECT 102.965 2030.000 131.065 2048.000 ;
        RECT 102.965 2029.000 105.000 2030.000 ;
      LAYER met4 ;
        RECT 0.000 2027.730 24.215 2029.000 ;
      LAYER met4 ;
        RECT 24.615 2027.330 104.600 2027.970 ;
      LAYER met4 ;
        RECT 105.000 2027.730 129.965 2030.000 ;
      LAYER met4 ;
        RECT 129.965 2029.000 131.065 2030.000 ;
        RECT 130.365 2027.330 131.065 2027.970 ;
      LAYER met4 ;
        RECT 131.465 2027.730 135.915 2559.270 ;
      LAYER met4 ;
        RECT 136.315 2558.965 136.915 2559.670 ;
        RECT 136.315 2029.000 136.915 2554.000 ;
        RECT 136.315 2027.330 136.915 2027.970 ;
      LAYER met4 ;
        RECT 137.315 2027.730 141.765 2559.270 ;
      LAYER met4 ;
        RECT 142.165 2558.965 142.865 2559.670 ;
        RECT 142.165 2029.000 142.865 2558.000 ;
        RECT 142.165 2027.330 142.865 2027.970 ;
        RECT 0.000 1995.690 142.865 2027.330 ;
      LAYER met4 ;
        RECT 143.265 1996.090 143.595 2560.610 ;
      LAYER met4 ;
        RECT 0.000 1987.360 143.495 1995.690 ;
      LAYER met4 ;
        RECT 143.895 1987.760 146.875 2594.440 ;
      LAYER met4 ;
        RECT 147.275 2559.670 148.255 2594.840 ;
      LAYER met4 ;
        RECT 147.175 2558.000 148.355 2559.270 ;
      LAYER met4 ;
        RECT 147.275 2029.000 148.255 2558.000 ;
      LAYER met4 ;
        RECT 147.175 2027.730 148.355 2029.000 ;
      LAYER met4 ;
        RECT 147.275 2003.065 148.255 2027.330 ;
      LAYER met4 ;
        RECT 148.655 2003.465 151.635 2610.145 ;
        RECT 151.935 2605.090 152.265 3169.610 ;
      LAYER met4 ;
        RECT 152.665 3168.670 199.465 3170.010 ;
        RECT 152.665 3167.965 153.365 3168.670 ;
        RECT 152.665 2636.330 153.365 2636.970 ;
      LAYER met4 ;
        RECT 153.765 2636.730 158.415 3168.270 ;
      LAYER met4 ;
        RECT 158.815 3167.965 159.415 3168.670 ;
        RECT 158.815 2636.330 159.415 2636.970 ;
      LAYER met4 ;
        RECT 159.815 2636.730 163.265 3168.270 ;
      LAYER met4 ;
        RECT 163.665 3167.965 164.265 3168.670 ;
        RECT 163.665 2636.330 164.265 2636.970 ;
      LAYER met4 ;
        RECT 164.665 2636.730 168.115 3168.270 ;
      LAYER met4 ;
        RECT 168.515 3167.965 169.115 3168.670 ;
        RECT 168.515 2636.330 169.115 2636.970 ;
      LAYER met4 ;
        RECT 169.515 2636.730 174.165 3168.270 ;
      LAYER met4 ;
        RECT 174.565 3167.965 175.165 3168.670 ;
        RECT 180.615 3168.365 186.065 3168.670 ;
        RECT 174.565 2636.330 175.165 2636.970 ;
      LAYER met4 ;
        RECT 175.565 2636.730 180.215 3168.270 ;
      LAYER met4 ;
        RECT 180.615 3167.965 181.215 3168.365 ;
        RECT 185.465 3167.965 186.065 3168.365 ;
      LAYER met4 ;
        RECT 181.615 2636.970 185.065 3167.965 ;
      LAYER met4 ;
        RECT 180.615 2636.570 181.215 2636.970 ;
        RECT 185.465 2636.570 186.065 2636.970 ;
      LAYER met4 ;
        RECT 186.465 2636.730 191.115 3168.270 ;
      LAYER met4 ;
        RECT 191.515 3167.965 192.115 3168.670 ;
        RECT 180.615 2636.330 186.065 2636.570 ;
        RECT 191.515 2636.330 192.115 2636.970 ;
      LAYER met4 ;
        RECT 192.515 2636.730 197.965 3168.270 ;
      LAYER met4 ;
        RECT 198.365 3167.965 199.465 3168.670 ;
      LAYER met4 ;
        RECT 3383.150 3140.050 3383.450 3214.550 ;
      LAYER met4 ;
        RECT 3388.535 3196.310 3435.965 3239.990 ;
        RECT 3388.535 3164.670 3435.335 3196.310 ;
        RECT 3388.535 3164.030 3389.635 3164.670 ;
      LAYER met4 ;
        RECT 3381.310 3139.750 3383.450 3140.050 ;
        RECT 3381.310 3021.050 3381.610 3139.750 ;
        RECT 3381.310 3020.750 3382.530 3021.050 ;
        RECT 3382.230 2898.650 3382.530 3020.750 ;
        RECT 3382.230 2898.350 3383.450 2898.650 ;
        RECT 3383.150 2800.050 3383.450 2898.350 ;
        RECT 3383.150 2799.750 3387.130 2800.050 ;
        RECT 3386.830 2732.490 3387.130 2799.750 ;
        RECT 3380.870 2731.310 3382.050 2732.490 ;
        RECT 3386.390 2731.310 3387.570 2732.490 ;
        RECT 3381.310 2705.290 3381.610 2731.310 ;
        RECT 3380.870 2704.110 3382.050 2705.290 ;
        RECT 3385.470 2704.110 3386.650 2705.290 ;
      LAYER met4 ;
        RECT 198.365 2636.330 199.465 2636.970 ;
        RECT 152.665 2604.690 199.465 2636.330 ;
      LAYER met4 ;
        RECT 3385.910 2609.650 3386.210 2704.110 ;
      LAYER met4 ;
        RECT 152.035 2561.010 199.465 2604.690 ;
        RECT 147.275 2001.545 151.535 2003.065 ;
        RECT 147.275 1987.360 148.255 2001.545 ;
        RECT 0.000 1985.840 148.255 1987.360 ;
        RECT 0.000 1952.010 143.495 1985.840 ;
        RECT 0.000 1950.670 142.865 1952.010 ;
      LAYER met4 ;
        RECT 0.000 1949.000 24.215 1950.270 ;
      LAYER met4 ;
        RECT 24.615 1949.965 104.600 1950.670 ;
        RECT 0.000 1421.000 25.965 1949.000 ;
        RECT 102.965 1945.000 105.000 1949.000 ;
      LAYER met4 ;
        RECT 105.000 1945.000 129.965 1950.270 ;
      LAYER met4 ;
        RECT 130.365 1949.965 131.065 1950.670 ;
        RECT 129.965 1945.000 131.065 1949.000 ;
        RECT 102.965 1942.000 131.065 1945.000 ;
        RECT 102.965 1940.000 105.000 1942.000 ;
      LAYER met4 ;
        RECT 105.000 1940.000 129.965 1942.000 ;
      LAYER met4 ;
        RECT 129.965 1940.000 131.065 1942.000 ;
        RECT 102.965 1922.000 131.065 1940.000 ;
        RECT 102.965 1920.000 105.000 1922.000 ;
      LAYER met4 ;
        RECT 105.000 1920.000 129.965 1922.000 ;
      LAYER met4 ;
        RECT 129.965 1920.000 131.065 1922.000 ;
        RECT 102.965 1902.000 131.065 1920.000 ;
        RECT 102.965 1900.000 105.000 1902.000 ;
      LAYER met4 ;
        RECT 105.000 1900.000 129.965 1902.000 ;
      LAYER met4 ;
        RECT 129.965 1900.000 131.065 1902.000 ;
        RECT 102.965 1882.000 131.065 1900.000 ;
        RECT 102.965 1880.000 105.000 1882.000 ;
      LAYER met4 ;
        RECT 105.000 1880.000 129.965 1882.000 ;
      LAYER met4 ;
        RECT 129.965 1880.000 131.065 1882.000 ;
        RECT 102.965 1862.000 131.065 1880.000 ;
        RECT 102.965 1860.000 105.000 1862.000 ;
      LAYER met4 ;
        RECT 105.000 1860.000 129.965 1862.000 ;
      LAYER met4 ;
        RECT 129.965 1860.000 131.065 1862.000 ;
        RECT 102.965 1842.000 131.065 1860.000 ;
        RECT 102.965 1840.000 105.000 1842.000 ;
      LAYER met4 ;
        RECT 105.000 1840.000 129.965 1842.000 ;
      LAYER met4 ;
        RECT 129.965 1840.000 131.065 1842.000 ;
        RECT 102.965 1822.000 131.065 1840.000 ;
        RECT 102.965 1820.000 105.000 1822.000 ;
      LAYER met4 ;
        RECT 105.000 1820.000 129.965 1822.000 ;
      LAYER met4 ;
        RECT 129.965 1820.000 131.065 1822.000 ;
        RECT 102.965 1802.000 131.065 1820.000 ;
        RECT 102.965 1800.000 105.000 1802.000 ;
      LAYER met4 ;
        RECT 105.000 1800.000 129.965 1802.000 ;
      LAYER met4 ;
        RECT 129.965 1800.000 131.065 1802.000 ;
        RECT 102.965 1782.000 131.065 1800.000 ;
        RECT 102.965 1780.000 105.000 1782.000 ;
      LAYER met4 ;
        RECT 105.000 1780.000 129.965 1782.000 ;
      LAYER met4 ;
        RECT 129.965 1780.000 131.065 1782.000 ;
        RECT 102.965 1762.000 131.065 1780.000 ;
        RECT 102.965 1760.000 105.000 1762.000 ;
      LAYER met4 ;
        RECT 105.000 1760.000 129.965 1762.000 ;
      LAYER met4 ;
        RECT 129.965 1760.000 131.065 1762.000 ;
        RECT 102.965 1742.000 131.065 1760.000 ;
        RECT 102.965 1740.000 105.000 1742.000 ;
      LAYER met4 ;
        RECT 105.000 1740.000 129.965 1742.000 ;
      LAYER met4 ;
        RECT 129.965 1740.000 131.065 1742.000 ;
        RECT 102.965 1722.000 131.065 1740.000 ;
        RECT 102.965 1720.000 105.000 1722.000 ;
      LAYER met4 ;
        RECT 105.000 1720.000 129.965 1722.000 ;
      LAYER met4 ;
        RECT 129.965 1720.000 131.065 1722.000 ;
        RECT 102.965 1702.000 131.065 1720.000 ;
        RECT 102.965 1700.000 105.000 1702.000 ;
      LAYER met4 ;
        RECT 105.000 1700.000 129.965 1702.000 ;
      LAYER met4 ;
        RECT 129.965 1700.000 131.065 1702.000 ;
        RECT 102.965 1682.000 131.065 1700.000 ;
        RECT 102.965 1680.000 105.000 1682.000 ;
      LAYER met4 ;
        RECT 105.000 1680.000 129.965 1682.000 ;
      LAYER met4 ;
        RECT 129.965 1680.000 131.065 1682.000 ;
        RECT 102.965 1662.000 131.065 1680.000 ;
        RECT 102.965 1660.000 105.000 1662.000 ;
      LAYER met4 ;
        RECT 105.000 1660.000 129.965 1662.000 ;
      LAYER met4 ;
        RECT 129.965 1660.000 131.065 1662.000 ;
        RECT 102.965 1642.000 131.065 1660.000 ;
        RECT 102.965 1640.000 105.000 1642.000 ;
      LAYER met4 ;
        RECT 105.000 1640.000 129.965 1642.000 ;
      LAYER met4 ;
        RECT 129.965 1640.000 131.065 1642.000 ;
        RECT 102.965 1622.000 131.065 1640.000 ;
        RECT 102.965 1620.000 105.000 1622.000 ;
      LAYER met4 ;
        RECT 105.000 1620.000 129.965 1622.000 ;
      LAYER met4 ;
        RECT 129.965 1620.000 131.065 1622.000 ;
        RECT 102.965 1602.000 131.065 1620.000 ;
        RECT 102.965 1600.000 105.000 1602.000 ;
      LAYER met4 ;
        RECT 105.000 1600.000 129.965 1602.000 ;
      LAYER met4 ;
        RECT 129.965 1600.000 131.065 1602.000 ;
        RECT 102.965 1582.000 131.065 1600.000 ;
        RECT 102.965 1580.000 105.000 1582.000 ;
      LAYER met4 ;
        RECT 105.000 1580.000 129.965 1582.000 ;
      LAYER met4 ;
        RECT 129.965 1580.000 131.065 1582.000 ;
        RECT 102.965 1562.000 131.065 1580.000 ;
        RECT 102.965 1560.000 105.000 1562.000 ;
      LAYER met4 ;
        RECT 105.000 1560.000 129.965 1562.000 ;
      LAYER met4 ;
        RECT 129.965 1560.000 131.065 1562.000 ;
        RECT 102.965 1542.000 131.065 1560.000 ;
        RECT 102.965 1540.000 105.000 1542.000 ;
      LAYER met4 ;
        RECT 105.000 1540.000 129.965 1542.000 ;
      LAYER met4 ;
        RECT 129.965 1540.000 131.065 1542.000 ;
        RECT 102.965 1522.000 131.065 1540.000 ;
        RECT 102.965 1520.000 105.000 1522.000 ;
      LAYER met4 ;
        RECT 105.000 1520.000 129.965 1522.000 ;
      LAYER met4 ;
        RECT 129.965 1520.000 131.065 1522.000 ;
        RECT 102.965 1502.000 131.065 1520.000 ;
        RECT 102.965 1500.000 105.000 1502.000 ;
      LAYER met4 ;
        RECT 105.000 1500.000 129.965 1502.000 ;
      LAYER met4 ;
        RECT 129.965 1500.000 131.065 1502.000 ;
        RECT 102.965 1482.000 131.065 1500.000 ;
        RECT 102.965 1480.000 105.000 1482.000 ;
      LAYER met4 ;
        RECT 105.000 1480.000 129.965 1482.000 ;
      LAYER met4 ;
        RECT 129.965 1480.000 131.065 1482.000 ;
        RECT 102.965 1462.000 131.065 1480.000 ;
        RECT 102.965 1460.000 105.000 1462.000 ;
      LAYER met4 ;
        RECT 105.000 1460.000 129.965 1462.000 ;
      LAYER met4 ;
        RECT 129.965 1460.000 131.065 1462.000 ;
        RECT 102.965 1442.000 131.065 1460.000 ;
        RECT 102.965 1440.000 105.000 1442.000 ;
      LAYER met4 ;
        RECT 105.000 1440.000 129.965 1442.000 ;
      LAYER met4 ;
        RECT 129.965 1440.000 131.065 1442.000 ;
        RECT 102.965 1422.000 131.065 1440.000 ;
        RECT 102.965 1421.000 105.000 1422.000 ;
      LAYER met4 ;
        RECT 0.000 1419.730 24.215 1421.000 ;
      LAYER met4 ;
        RECT 24.615 1419.330 104.600 1419.970 ;
      LAYER met4 ;
        RECT 105.000 1419.730 129.965 1422.000 ;
      LAYER met4 ;
        RECT 129.965 1421.000 131.065 1422.000 ;
        RECT 130.365 1419.330 131.065 1419.970 ;
      LAYER met4 ;
        RECT 131.465 1419.730 135.915 1950.270 ;
      LAYER met4 ;
        RECT 136.315 1949.965 136.915 1950.670 ;
        RECT 136.315 1421.000 136.915 1946.000 ;
        RECT 136.315 1419.330 136.915 1419.970 ;
      LAYER met4 ;
        RECT 137.315 1419.730 141.765 1950.270 ;
      LAYER met4 ;
        RECT 142.165 1949.965 142.865 1950.670 ;
        RECT 142.165 1421.000 142.865 1949.000 ;
        RECT 142.165 1419.330 142.865 1419.970 ;
        RECT 0.000 1387.690 142.865 1419.330 ;
      LAYER met4 ;
        RECT 143.265 1388.090 143.595 1951.610 ;
      LAYER met4 ;
        RECT 0.000 1379.360 143.495 1387.690 ;
      LAYER met4 ;
        RECT 143.895 1379.760 146.875 1985.440 ;
      LAYER met4 ;
        RECT 147.275 1950.670 148.255 1985.840 ;
      LAYER met4 ;
        RECT 147.175 1949.000 148.355 1950.270 ;
      LAYER met4 ;
        RECT 147.275 1421.000 148.255 1949.000 ;
      LAYER met4 ;
        RECT 147.175 1419.730 148.355 1421.000 ;
      LAYER met4 ;
        RECT 147.275 1395.065 148.255 1419.330 ;
      LAYER met4 ;
        RECT 148.655 1395.465 151.635 2001.145 ;
        RECT 151.935 1996.090 152.265 2560.610 ;
      LAYER met4 ;
        RECT 152.665 2559.670 199.465 2561.010 ;
        RECT 152.665 2558.965 153.365 2559.670 ;
        RECT 152.665 2027.330 153.365 2027.970 ;
      LAYER met4 ;
        RECT 153.765 2027.730 158.415 2559.270 ;
      LAYER met4 ;
        RECT 158.815 2558.965 159.415 2559.670 ;
        RECT 158.815 2027.330 159.415 2027.970 ;
      LAYER met4 ;
        RECT 159.815 2027.730 163.265 2559.270 ;
      LAYER met4 ;
        RECT 163.665 2558.965 164.265 2559.670 ;
        RECT 163.665 2027.330 164.265 2027.970 ;
      LAYER met4 ;
        RECT 164.665 2027.730 168.115 2559.270 ;
      LAYER met4 ;
        RECT 168.515 2558.965 169.115 2559.670 ;
        RECT 168.515 2027.330 169.115 2027.970 ;
      LAYER met4 ;
        RECT 169.515 2027.730 174.165 2559.270 ;
      LAYER met4 ;
        RECT 174.565 2558.965 175.165 2559.670 ;
        RECT 180.615 2559.365 186.065 2559.670 ;
        RECT 174.565 2027.330 175.165 2027.970 ;
      LAYER met4 ;
        RECT 175.565 2027.730 180.215 2559.270 ;
      LAYER met4 ;
        RECT 180.615 2558.965 181.215 2559.365 ;
        RECT 185.465 2558.965 186.065 2559.365 ;
      LAYER met4 ;
        RECT 181.615 2027.970 185.065 2558.965 ;
      LAYER met4 ;
        RECT 180.615 2027.570 181.215 2027.970 ;
        RECT 185.465 2027.570 186.065 2027.970 ;
      LAYER met4 ;
        RECT 186.465 2027.730 191.115 2559.270 ;
      LAYER met4 ;
        RECT 191.515 2558.965 192.115 2559.670 ;
        RECT 180.615 2027.330 186.065 2027.570 ;
        RECT 191.515 2027.330 192.115 2027.970 ;
      LAYER met4 ;
        RECT 192.515 2027.730 197.965 2559.270 ;
      LAYER met4 ;
        RECT 198.365 2558.965 199.465 2559.670 ;
      LAYER met4 ;
        RECT 3383.150 2609.350 3386.210 2609.650 ;
      LAYER met4 ;
        RECT 3388.535 2632.330 3389.635 2633.035 ;
      LAYER met4 ;
        RECT 3390.035 2632.730 3395.485 3164.270 ;
      LAYER met4 ;
        RECT 3395.885 3164.030 3396.485 3164.670 ;
        RECT 3401.935 3164.430 3407.385 3164.670 ;
        RECT 3395.885 2632.330 3396.485 2633.035 ;
      LAYER met4 ;
        RECT 3396.885 2632.730 3401.535 3164.270 ;
      LAYER met4 ;
        RECT 3401.935 3164.030 3402.535 3164.430 ;
        RECT 3406.785 3164.030 3407.385 3164.430 ;
      LAYER met4 ;
        RECT 3402.935 2633.035 3406.385 3164.030 ;
      LAYER met4 ;
        RECT 3401.935 2632.635 3402.535 2633.035 ;
        RECT 3406.785 2632.635 3407.385 2633.035 ;
      LAYER met4 ;
        RECT 3407.785 2632.730 3412.435 3164.270 ;
      LAYER met4 ;
        RECT 3412.835 3164.030 3413.435 3164.670 ;
        RECT 3401.935 2632.330 3407.385 2632.635 ;
        RECT 3412.835 2632.330 3413.435 2633.035 ;
      LAYER met4 ;
        RECT 3413.835 2632.730 3418.485 3164.270 ;
      LAYER met4 ;
        RECT 3418.885 3164.030 3419.485 3164.670 ;
        RECT 3418.885 2632.330 3419.485 2633.035 ;
      LAYER met4 ;
        RECT 3419.885 2632.730 3423.335 3164.270 ;
      LAYER met4 ;
        RECT 3423.735 3164.030 3424.335 3164.670 ;
        RECT 3423.735 2632.330 3424.335 2633.035 ;
      LAYER met4 ;
        RECT 3424.735 2632.730 3428.185 3164.270 ;
      LAYER met4 ;
        RECT 3428.585 3164.030 3429.185 3164.670 ;
        RECT 3428.585 2632.330 3429.185 2633.035 ;
      LAYER met4 ;
        RECT 3429.585 2632.730 3434.235 3164.270 ;
      LAYER met4 ;
        RECT 3434.635 3164.030 3435.335 3164.670 ;
        RECT 3434.635 2632.330 3435.335 2633.035 ;
        RECT 3388.535 2630.990 3435.335 2632.330 ;
      LAYER met4 ;
        RECT 3435.735 2631.390 3436.065 3195.910 ;
        RECT 3436.365 3190.855 3439.345 3796.535 ;
      LAYER met4 ;
        RECT 3439.745 3772.670 3440.725 3796.935 ;
      LAYER met4 ;
        RECT 3439.645 3771.000 3440.825 3772.270 ;
      LAYER met4 ;
        RECT 3439.745 3243.000 3440.725 3771.000 ;
      LAYER met4 ;
        RECT 3439.645 3241.730 3440.825 3243.000 ;
      LAYER met4 ;
        RECT 3439.745 3206.160 3440.725 3241.330 ;
      LAYER met4 ;
        RECT 3441.125 3206.560 3444.105 3812.240 ;
      LAYER met4 ;
        RECT 3444.505 3804.310 3588.000 3812.640 ;
      LAYER met4 ;
        RECT 3444.405 3240.390 3444.735 3803.910 ;
      LAYER met4 ;
        RECT 3445.135 3772.670 3588.000 3804.310 ;
        RECT 3445.135 3772.030 3445.835 3772.670 ;
        RECT 3445.135 3243.000 3445.835 3771.000 ;
        RECT 3445.135 3241.330 3445.835 3242.035 ;
      LAYER met4 ;
        RECT 3446.235 3241.730 3450.685 3772.270 ;
      LAYER met4 ;
        RECT 3451.085 3772.030 3451.685 3772.670 ;
        RECT 3451.085 3243.000 3451.685 3768.000 ;
        RECT 3451.085 3241.330 3451.685 3242.035 ;
      LAYER met4 ;
        RECT 3452.085 3241.730 3456.535 3772.270 ;
      LAYER met4 ;
        RECT 3456.935 3772.030 3457.635 3772.670 ;
        RECT 3456.935 3767.000 3458.035 3771.000 ;
      LAYER met4 ;
        RECT 3458.035 3767.000 3483.000 3772.270 ;
      LAYER met4 ;
        RECT 3483.400 3772.030 3563.385 3772.670 ;
      LAYER met4 ;
        RECT 3563.785 3771.000 3588.000 3772.270 ;
      LAYER met4 ;
        RECT 3483.000 3767.000 3485.035 3771.000 ;
        RECT 3456.935 3764.000 3485.035 3767.000 ;
        RECT 3456.935 3762.000 3458.035 3764.000 ;
      LAYER met4 ;
        RECT 3458.035 3762.000 3483.000 3764.000 ;
      LAYER met4 ;
        RECT 3483.000 3762.000 3485.035 3764.000 ;
        RECT 3456.935 3744.000 3485.035 3762.000 ;
        RECT 3456.935 3742.000 3458.035 3744.000 ;
      LAYER met4 ;
        RECT 3458.035 3742.000 3483.000 3744.000 ;
      LAYER met4 ;
        RECT 3483.000 3742.000 3485.035 3744.000 ;
        RECT 3456.935 3724.000 3485.035 3742.000 ;
        RECT 3456.935 3722.000 3458.035 3724.000 ;
      LAYER met4 ;
        RECT 3458.035 3722.000 3483.000 3724.000 ;
      LAYER met4 ;
        RECT 3483.000 3722.000 3485.035 3724.000 ;
        RECT 3456.935 3704.000 3485.035 3722.000 ;
        RECT 3456.935 3702.000 3458.035 3704.000 ;
      LAYER met4 ;
        RECT 3458.035 3702.000 3483.000 3704.000 ;
      LAYER met4 ;
        RECT 3483.000 3702.000 3485.035 3704.000 ;
        RECT 3456.935 3684.000 3485.035 3702.000 ;
        RECT 3456.935 3682.000 3458.035 3684.000 ;
      LAYER met4 ;
        RECT 3458.035 3682.000 3483.000 3684.000 ;
      LAYER met4 ;
        RECT 3483.000 3682.000 3485.035 3684.000 ;
        RECT 3456.935 3664.000 3485.035 3682.000 ;
        RECT 3456.935 3662.000 3458.035 3664.000 ;
      LAYER met4 ;
        RECT 3458.035 3662.000 3483.000 3664.000 ;
      LAYER met4 ;
        RECT 3483.000 3662.000 3485.035 3664.000 ;
        RECT 3456.935 3644.000 3485.035 3662.000 ;
        RECT 3456.935 3642.000 3458.035 3644.000 ;
      LAYER met4 ;
        RECT 3458.035 3642.000 3483.000 3644.000 ;
      LAYER met4 ;
        RECT 3483.000 3642.000 3485.035 3644.000 ;
        RECT 3456.935 3624.000 3485.035 3642.000 ;
        RECT 3456.935 3622.000 3458.035 3624.000 ;
      LAYER met4 ;
        RECT 3458.035 3622.000 3483.000 3624.000 ;
      LAYER met4 ;
        RECT 3483.000 3622.000 3485.035 3624.000 ;
        RECT 3456.935 3604.000 3485.035 3622.000 ;
        RECT 3456.935 3602.000 3458.035 3604.000 ;
      LAYER met4 ;
        RECT 3458.035 3602.000 3483.000 3604.000 ;
      LAYER met4 ;
        RECT 3483.000 3602.000 3485.035 3604.000 ;
        RECT 3456.935 3584.000 3485.035 3602.000 ;
        RECT 3456.935 3582.000 3458.035 3584.000 ;
      LAYER met4 ;
        RECT 3458.035 3582.000 3483.000 3584.000 ;
      LAYER met4 ;
        RECT 3483.000 3582.000 3485.035 3584.000 ;
        RECT 3456.935 3564.000 3485.035 3582.000 ;
        RECT 3456.935 3562.000 3458.035 3564.000 ;
      LAYER met4 ;
        RECT 3458.035 3562.000 3483.000 3564.000 ;
      LAYER met4 ;
        RECT 3483.000 3562.000 3485.035 3564.000 ;
        RECT 3456.935 3544.000 3485.035 3562.000 ;
        RECT 3456.935 3542.000 3458.035 3544.000 ;
      LAYER met4 ;
        RECT 3458.035 3542.000 3483.000 3544.000 ;
      LAYER met4 ;
        RECT 3483.000 3542.000 3485.035 3544.000 ;
        RECT 3456.935 3524.000 3485.035 3542.000 ;
        RECT 3456.935 3522.000 3458.035 3524.000 ;
      LAYER met4 ;
        RECT 3458.035 3522.000 3483.000 3524.000 ;
      LAYER met4 ;
        RECT 3483.000 3522.000 3485.035 3524.000 ;
        RECT 3456.935 3504.000 3485.035 3522.000 ;
        RECT 3456.935 3502.000 3458.035 3504.000 ;
      LAYER met4 ;
        RECT 3458.035 3502.000 3483.000 3504.000 ;
      LAYER met4 ;
        RECT 3483.000 3502.000 3485.035 3504.000 ;
        RECT 3456.935 3484.000 3485.035 3502.000 ;
        RECT 3456.935 3482.000 3458.035 3484.000 ;
      LAYER met4 ;
        RECT 3458.035 3482.000 3483.000 3484.000 ;
      LAYER met4 ;
        RECT 3483.000 3482.000 3485.035 3484.000 ;
        RECT 3456.935 3464.000 3485.035 3482.000 ;
        RECT 3456.935 3462.000 3458.035 3464.000 ;
      LAYER met4 ;
        RECT 3458.035 3462.000 3483.000 3464.000 ;
      LAYER met4 ;
        RECT 3483.000 3462.000 3485.035 3464.000 ;
        RECT 3456.935 3444.000 3485.035 3462.000 ;
        RECT 3456.935 3442.000 3458.035 3444.000 ;
      LAYER met4 ;
        RECT 3458.035 3442.000 3483.000 3444.000 ;
      LAYER met4 ;
        RECT 3483.000 3442.000 3485.035 3444.000 ;
        RECT 3456.935 3424.000 3485.035 3442.000 ;
        RECT 3456.935 3422.000 3458.035 3424.000 ;
      LAYER met4 ;
        RECT 3458.035 3422.000 3483.000 3424.000 ;
      LAYER met4 ;
        RECT 3483.000 3422.000 3485.035 3424.000 ;
        RECT 3456.935 3404.000 3485.035 3422.000 ;
        RECT 3456.935 3402.000 3458.035 3404.000 ;
      LAYER met4 ;
        RECT 3458.035 3402.000 3483.000 3404.000 ;
      LAYER met4 ;
        RECT 3483.000 3402.000 3485.035 3404.000 ;
        RECT 3456.935 3384.000 3485.035 3402.000 ;
        RECT 3456.935 3382.000 3458.035 3384.000 ;
      LAYER met4 ;
        RECT 3458.035 3382.000 3483.000 3384.000 ;
      LAYER met4 ;
        RECT 3483.000 3382.000 3485.035 3384.000 ;
        RECT 3456.935 3364.000 3485.035 3382.000 ;
        RECT 3456.935 3362.000 3458.035 3364.000 ;
      LAYER met4 ;
        RECT 3458.035 3362.000 3483.000 3364.000 ;
      LAYER met4 ;
        RECT 3483.000 3362.000 3485.035 3364.000 ;
        RECT 3456.935 3344.000 3485.035 3362.000 ;
        RECT 3456.935 3342.000 3458.035 3344.000 ;
      LAYER met4 ;
        RECT 3458.035 3342.000 3483.000 3344.000 ;
      LAYER met4 ;
        RECT 3483.000 3342.000 3485.035 3344.000 ;
        RECT 3456.935 3324.000 3485.035 3342.000 ;
        RECT 3456.935 3322.000 3458.035 3324.000 ;
      LAYER met4 ;
        RECT 3458.035 3322.000 3483.000 3324.000 ;
      LAYER met4 ;
        RECT 3483.000 3322.000 3485.035 3324.000 ;
        RECT 3456.935 3304.000 3485.035 3322.000 ;
        RECT 3456.935 3302.000 3458.035 3304.000 ;
      LAYER met4 ;
        RECT 3458.035 3302.000 3483.000 3304.000 ;
      LAYER met4 ;
        RECT 3483.000 3302.000 3485.035 3304.000 ;
        RECT 3456.935 3284.000 3485.035 3302.000 ;
        RECT 3456.935 3282.000 3458.035 3284.000 ;
      LAYER met4 ;
        RECT 3458.035 3282.000 3483.000 3284.000 ;
      LAYER met4 ;
        RECT 3483.000 3282.000 3485.035 3284.000 ;
        RECT 3456.935 3264.000 3485.035 3282.000 ;
        RECT 3456.935 3262.000 3458.035 3264.000 ;
      LAYER met4 ;
        RECT 3458.035 3262.000 3483.000 3264.000 ;
      LAYER met4 ;
        RECT 3483.000 3262.000 3485.035 3264.000 ;
        RECT 3456.935 3244.000 3485.035 3262.000 ;
        RECT 3456.935 3243.000 3458.035 3244.000 ;
        RECT 3456.935 3241.330 3457.635 3242.035 ;
      LAYER met4 ;
        RECT 3458.035 3241.730 3483.000 3244.000 ;
      LAYER met4 ;
        RECT 3483.000 3243.000 3485.035 3244.000 ;
        RECT 3562.035 3243.000 3588.000 3771.000 ;
        RECT 3483.400 3241.330 3563.385 3242.035 ;
      LAYER met4 ;
        RECT 3563.785 3241.730 3588.000 3243.000 ;
      LAYER met4 ;
        RECT 3445.135 3239.990 3588.000 3241.330 ;
        RECT 3444.505 3206.160 3588.000 3239.990 ;
        RECT 3439.745 3204.640 3588.000 3206.160 ;
        RECT 3439.745 3190.455 3440.725 3204.640 ;
        RECT 3436.465 3188.935 3440.725 3190.455 ;
      LAYER met4 ;
        RECT 3383.150 2555.250 3383.450 2609.350 ;
        RECT 3382.230 2554.950 3383.450 2555.250 ;
      LAYER met4 ;
        RECT 3388.535 2587.310 3435.965 2630.990 ;
        RECT 3388.535 2555.670 3435.335 2587.310 ;
        RECT 3388.535 2555.030 3389.635 2555.670 ;
      LAYER met4 ;
        RECT 3382.230 2511.050 3382.530 2554.950 ;
        RECT 3382.230 2510.750 3383.450 2511.050 ;
        RECT 3383.150 2415.850 3383.450 2510.750 ;
        RECT 3383.150 2415.550 3386.210 2415.850 ;
        RECT 3385.910 2344.450 3386.210 2415.550 ;
        RECT 3384.990 2344.150 3386.210 2344.450 ;
        RECT 3384.990 2249.250 3385.290 2344.150 ;
        RECT 3382.230 2248.950 3385.290 2249.250 ;
        RECT 3382.230 2150.650 3382.530 2248.950 ;
        RECT 3381.310 2150.350 3382.530 2150.650 ;
        RECT 3381.310 2055.450 3381.610 2150.350 ;
        RECT 3381.310 2055.150 3383.450 2055.450 ;
      LAYER met4 ;
        RECT 198.365 2027.330 199.465 2027.970 ;
        RECT 152.665 1995.690 199.465 2027.330 ;
        RECT 152.035 1952.010 199.465 1995.690 ;
      LAYER met4 ;
        RECT 3369.335 1958.575 3369.665 1958.905 ;
      LAYER met4 ;
        RECT 147.275 1393.545 151.535 1395.065 ;
        RECT 147.275 1379.360 148.255 1393.545 ;
        RECT 0.000 1377.840 148.255 1379.360 ;
        RECT 0.000 1344.010 143.495 1377.840 ;
        RECT 0.000 1342.670 142.865 1344.010 ;
      LAYER met4 ;
        RECT 0.000 1341.000 24.215 1342.270 ;
      LAYER met4 ;
        RECT 24.615 1341.965 104.600 1342.670 ;
        RECT 0.000 812.000 25.965 1341.000 ;
        RECT 102.965 1336.000 105.000 1341.000 ;
      LAYER met4 ;
        RECT 105.000 1336.000 129.965 1342.270 ;
      LAYER met4 ;
        RECT 130.365 1341.965 131.065 1342.670 ;
        RECT 129.965 1336.000 131.065 1341.000 ;
        RECT 102.965 1333.000 131.065 1336.000 ;
        RECT 102.965 1331.000 105.000 1333.000 ;
      LAYER met4 ;
        RECT 105.000 1331.000 129.965 1333.000 ;
      LAYER met4 ;
        RECT 129.965 1331.000 131.065 1333.000 ;
        RECT 102.965 1313.000 131.065 1331.000 ;
        RECT 102.965 1311.000 105.000 1313.000 ;
      LAYER met4 ;
        RECT 105.000 1311.000 129.965 1313.000 ;
      LAYER met4 ;
        RECT 129.965 1311.000 131.065 1313.000 ;
        RECT 102.965 1293.000 131.065 1311.000 ;
        RECT 102.965 1291.000 105.000 1293.000 ;
      LAYER met4 ;
        RECT 105.000 1291.000 129.965 1293.000 ;
      LAYER met4 ;
        RECT 129.965 1291.000 131.065 1293.000 ;
        RECT 102.965 1273.000 131.065 1291.000 ;
        RECT 102.965 1271.000 105.000 1273.000 ;
      LAYER met4 ;
        RECT 105.000 1271.000 129.965 1273.000 ;
      LAYER met4 ;
        RECT 129.965 1271.000 131.065 1273.000 ;
        RECT 102.965 1253.000 131.065 1271.000 ;
        RECT 102.965 1251.000 105.000 1253.000 ;
      LAYER met4 ;
        RECT 105.000 1251.000 129.965 1253.000 ;
      LAYER met4 ;
        RECT 129.965 1251.000 131.065 1253.000 ;
        RECT 102.965 1233.000 131.065 1251.000 ;
        RECT 102.965 1231.000 105.000 1233.000 ;
      LAYER met4 ;
        RECT 105.000 1231.000 129.965 1233.000 ;
      LAYER met4 ;
        RECT 129.965 1231.000 131.065 1233.000 ;
        RECT 102.965 1213.000 131.065 1231.000 ;
        RECT 102.965 1211.000 105.000 1213.000 ;
      LAYER met4 ;
        RECT 105.000 1211.000 129.965 1213.000 ;
      LAYER met4 ;
        RECT 129.965 1211.000 131.065 1213.000 ;
        RECT 102.965 1193.000 131.065 1211.000 ;
        RECT 102.965 1191.000 105.000 1193.000 ;
      LAYER met4 ;
        RECT 105.000 1191.000 129.965 1193.000 ;
      LAYER met4 ;
        RECT 129.965 1191.000 131.065 1193.000 ;
        RECT 102.965 1173.000 131.065 1191.000 ;
        RECT 102.965 1171.000 105.000 1173.000 ;
      LAYER met4 ;
        RECT 105.000 1171.000 129.965 1173.000 ;
      LAYER met4 ;
        RECT 129.965 1171.000 131.065 1173.000 ;
        RECT 102.965 1153.000 131.065 1171.000 ;
        RECT 102.965 1151.000 105.000 1153.000 ;
      LAYER met4 ;
        RECT 105.000 1151.000 129.965 1153.000 ;
      LAYER met4 ;
        RECT 129.965 1151.000 131.065 1153.000 ;
        RECT 102.965 1133.000 131.065 1151.000 ;
        RECT 102.965 1131.000 105.000 1133.000 ;
      LAYER met4 ;
        RECT 105.000 1131.000 129.965 1133.000 ;
      LAYER met4 ;
        RECT 129.965 1131.000 131.065 1133.000 ;
        RECT 102.965 1113.000 131.065 1131.000 ;
        RECT 102.965 1111.000 105.000 1113.000 ;
      LAYER met4 ;
        RECT 105.000 1111.000 129.965 1113.000 ;
      LAYER met4 ;
        RECT 129.965 1111.000 131.065 1113.000 ;
        RECT 102.965 1093.000 131.065 1111.000 ;
        RECT 102.965 1091.000 105.000 1093.000 ;
      LAYER met4 ;
        RECT 105.000 1091.000 129.965 1093.000 ;
      LAYER met4 ;
        RECT 129.965 1091.000 131.065 1093.000 ;
        RECT 102.965 1073.000 131.065 1091.000 ;
        RECT 102.965 1071.000 105.000 1073.000 ;
      LAYER met4 ;
        RECT 105.000 1071.000 129.965 1073.000 ;
      LAYER met4 ;
        RECT 129.965 1071.000 131.065 1073.000 ;
        RECT 102.965 1053.000 131.065 1071.000 ;
        RECT 102.965 1051.000 105.000 1053.000 ;
      LAYER met4 ;
        RECT 105.000 1051.000 129.965 1053.000 ;
      LAYER met4 ;
        RECT 129.965 1051.000 131.065 1053.000 ;
        RECT 102.965 1033.000 131.065 1051.000 ;
        RECT 102.965 1031.000 105.000 1033.000 ;
      LAYER met4 ;
        RECT 105.000 1031.000 129.965 1033.000 ;
      LAYER met4 ;
        RECT 129.965 1031.000 131.065 1033.000 ;
        RECT 102.965 1013.000 131.065 1031.000 ;
        RECT 102.965 1011.000 105.000 1013.000 ;
      LAYER met4 ;
        RECT 105.000 1011.000 129.965 1013.000 ;
      LAYER met4 ;
        RECT 129.965 1011.000 131.065 1013.000 ;
        RECT 102.965 993.000 131.065 1011.000 ;
        RECT 102.965 991.000 105.000 993.000 ;
      LAYER met4 ;
        RECT 105.000 991.000 129.965 993.000 ;
      LAYER met4 ;
        RECT 129.965 991.000 131.065 993.000 ;
        RECT 102.965 973.000 131.065 991.000 ;
        RECT 102.965 971.000 105.000 973.000 ;
      LAYER met4 ;
        RECT 105.000 971.000 129.965 973.000 ;
      LAYER met4 ;
        RECT 129.965 971.000 131.065 973.000 ;
        RECT 102.965 953.000 131.065 971.000 ;
        RECT 102.965 951.000 105.000 953.000 ;
      LAYER met4 ;
        RECT 105.000 951.000 129.965 953.000 ;
      LAYER met4 ;
        RECT 129.965 951.000 131.065 953.000 ;
        RECT 102.965 933.000 131.065 951.000 ;
        RECT 102.965 931.000 105.000 933.000 ;
      LAYER met4 ;
        RECT 105.000 931.000 129.965 933.000 ;
      LAYER met4 ;
        RECT 129.965 931.000 131.065 933.000 ;
        RECT 102.965 913.000 131.065 931.000 ;
        RECT 102.965 911.000 105.000 913.000 ;
      LAYER met4 ;
        RECT 105.000 911.000 129.965 913.000 ;
      LAYER met4 ;
        RECT 129.965 911.000 131.065 913.000 ;
        RECT 102.965 893.000 131.065 911.000 ;
        RECT 102.965 891.000 105.000 893.000 ;
      LAYER met4 ;
        RECT 105.000 891.000 129.965 893.000 ;
      LAYER met4 ;
        RECT 129.965 891.000 131.065 893.000 ;
        RECT 102.965 873.000 131.065 891.000 ;
        RECT 102.965 871.000 105.000 873.000 ;
      LAYER met4 ;
        RECT 105.000 871.000 129.965 873.000 ;
      LAYER met4 ;
        RECT 129.965 871.000 131.065 873.000 ;
        RECT 102.965 853.000 131.065 871.000 ;
        RECT 102.965 851.000 105.000 853.000 ;
      LAYER met4 ;
        RECT 105.000 851.000 129.965 853.000 ;
      LAYER met4 ;
        RECT 129.965 851.000 131.065 853.000 ;
        RECT 102.965 833.000 131.065 851.000 ;
        RECT 102.965 831.000 105.000 833.000 ;
      LAYER met4 ;
        RECT 105.000 831.000 129.965 833.000 ;
      LAYER met4 ;
        RECT 129.965 831.000 131.065 833.000 ;
        RECT 102.965 813.000 131.065 831.000 ;
        RECT 102.965 812.000 105.000 813.000 ;
      LAYER met4 ;
        RECT 0.000 810.730 24.215 812.000 ;
      LAYER met4 ;
        RECT 24.615 810.330 104.600 810.970 ;
      LAYER met4 ;
        RECT 105.000 810.730 129.965 813.000 ;
      LAYER met4 ;
        RECT 129.965 812.000 131.065 813.000 ;
        RECT 130.365 810.330 131.065 810.970 ;
      LAYER met4 ;
        RECT 131.465 810.730 135.915 1342.270 ;
      LAYER met4 ;
        RECT 136.315 1341.965 136.915 1342.670 ;
        RECT 136.315 812.000 136.915 1337.000 ;
        RECT 136.315 810.330 136.915 810.970 ;
      LAYER met4 ;
        RECT 137.315 810.730 141.765 1342.270 ;
      LAYER met4 ;
        RECT 142.165 1341.965 142.865 1342.670 ;
        RECT 142.165 812.000 142.865 1341.000 ;
        RECT 142.165 810.330 142.865 810.970 ;
        RECT 0.000 778.690 142.865 810.330 ;
      LAYER met4 ;
        RECT 143.265 779.090 143.595 1343.610 ;
      LAYER met4 ;
        RECT 0.000 770.360 143.495 778.690 ;
      LAYER met4 ;
        RECT 143.895 770.760 146.875 1377.440 ;
      LAYER met4 ;
        RECT 147.275 1342.670 148.255 1377.840 ;
      LAYER met4 ;
        RECT 147.175 1341.000 148.355 1342.270 ;
      LAYER met4 ;
        RECT 147.275 812.000 148.255 1341.000 ;
      LAYER met4 ;
        RECT 147.175 810.730 148.355 812.000 ;
      LAYER met4 ;
        RECT 147.275 786.065 148.255 810.330 ;
      LAYER met4 ;
        RECT 148.655 786.465 151.635 1393.145 ;
        RECT 151.935 1388.090 152.265 1951.610 ;
      LAYER met4 ;
        RECT 152.665 1950.670 199.465 1952.010 ;
        RECT 152.665 1949.965 153.365 1950.670 ;
        RECT 152.665 1419.330 153.365 1419.970 ;
      LAYER met4 ;
        RECT 153.765 1419.730 158.415 1950.270 ;
      LAYER met4 ;
        RECT 158.815 1949.965 159.415 1950.670 ;
        RECT 158.815 1419.330 159.415 1419.970 ;
      LAYER met4 ;
        RECT 159.815 1419.730 163.265 1950.270 ;
      LAYER met4 ;
        RECT 163.665 1949.965 164.265 1950.670 ;
        RECT 163.665 1419.330 164.265 1419.970 ;
      LAYER met4 ;
        RECT 164.665 1419.730 168.115 1950.270 ;
      LAYER met4 ;
        RECT 168.515 1949.965 169.115 1950.670 ;
        RECT 168.515 1419.330 169.115 1419.970 ;
      LAYER met4 ;
        RECT 169.515 1419.730 174.165 1950.270 ;
      LAYER met4 ;
        RECT 174.565 1949.965 175.165 1950.670 ;
        RECT 180.615 1950.365 186.065 1950.670 ;
        RECT 174.565 1419.330 175.165 1419.970 ;
      LAYER met4 ;
        RECT 175.565 1419.730 180.215 1950.270 ;
      LAYER met4 ;
        RECT 180.615 1949.965 181.215 1950.365 ;
        RECT 185.465 1949.965 186.065 1950.365 ;
      LAYER met4 ;
        RECT 181.615 1419.970 185.065 1949.965 ;
      LAYER met4 ;
        RECT 180.615 1419.570 181.215 1419.970 ;
        RECT 185.465 1419.570 186.065 1419.970 ;
      LAYER met4 ;
        RECT 186.465 1419.730 191.115 1950.270 ;
      LAYER met4 ;
        RECT 191.515 1949.965 192.115 1950.670 ;
        RECT 180.615 1419.330 186.065 1419.570 ;
        RECT 191.515 1419.330 192.115 1419.970 ;
      LAYER met4 ;
        RECT 192.515 1419.730 197.965 1950.270 ;
      LAYER met4 ;
        RECT 198.365 1949.965 199.465 1950.670 ;
      LAYER met4 ;
        RECT 3369.350 1932.385 3369.650 1958.575 ;
        RECT 3383.150 1956.850 3383.450 2055.150 ;
        RECT 3382.230 1956.550 3383.450 1956.850 ;
      LAYER met4 ;
        RECT 3388.535 2023.330 3389.635 2024.035 ;
      LAYER met4 ;
        RECT 3390.035 2023.730 3395.485 2555.270 ;
      LAYER met4 ;
        RECT 3395.885 2555.030 3396.485 2555.670 ;
        RECT 3401.935 2555.430 3407.385 2555.670 ;
        RECT 3395.885 2023.330 3396.485 2024.035 ;
      LAYER met4 ;
        RECT 3396.885 2023.730 3401.535 2555.270 ;
      LAYER met4 ;
        RECT 3401.935 2555.030 3402.535 2555.430 ;
        RECT 3406.785 2555.030 3407.385 2555.430 ;
      LAYER met4 ;
        RECT 3402.935 2024.035 3406.385 2555.030 ;
      LAYER met4 ;
        RECT 3401.935 2023.635 3402.535 2024.035 ;
        RECT 3406.785 2023.635 3407.385 2024.035 ;
      LAYER met4 ;
        RECT 3407.785 2023.730 3412.435 2555.270 ;
      LAYER met4 ;
        RECT 3412.835 2555.030 3413.435 2555.670 ;
        RECT 3401.935 2023.330 3407.385 2023.635 ;
        RECT 3412.835 2023.330 3413.435 2024.035 ;
      LAYER met4 ;
        RECT 3413.835 2023.730 3418.485 2555.270 ;
      LAYER met4 ;
        RECT 3418.885 2555.030 3419.485 2555.670 ;
        RECT 3418.885 2023.330 3419.485 2024.035 ;
      LAYER met4 ;
        RECT 3419.885 2023.730 3423.335 2555.270 ;
      LAYER met4 ;
        RECT 3423.735 2555.030 3424.335 2555.670 ;
        RECT 3423.735 2023.330 3424.335 2024.035 ;
      LAYER met4 ;
        RECT 3424.735 2023.730 3428.185 2555.270 ;
      LAYER met4 ;
        RECT 3428.585 2555.030 3429.185 2555.670 ;
        RECT 3428.585 2023.330 3429.185 2024.035 ;
      LAYER met4 ;
        RECT 3429.585 2023.730 3434.235 2555.270 ;
      LAYER met4 ;
        RECT 3434.635 2555.030 3435.335 2555.670 ;
        RECT 3434.635 2023.330 3435.335 2024.035 ;
        RECT 3388.535 2021.990 3435.335 2023.330 ;
      LAYER met4 ;
        RECT 3435.735 2022.390 3436.065 2586.910 ;
        RECT 3436.365 2581.855 3439.345 3188.535 ;
      LAYER met4 ;
        RECT 3439.745 3164.670 3440.725 3188.935 ;
      LAYER met4 ;
        RECT 3439.645 3163.000 3440.825 3164.270 ;
      LAYER met4 ;
        RECT 3439.745 2634.000 3440.725 3163.000 ;
      LAYER met4 ;
        RECT 3439.645 2632.730 3440.825 2634.000 ;
      LAYER met4 ;
        RECT 3439.745 2597.160 3440.725 2632.330 ;
      LAYER met4 ;
        RECT 3441.125 2597.560 3444.105 3204.240 ;
      LAYER met4 ;
        RECT 3444.505 3196.310 3588.000 3204.640 ;
      LAYER met4 ;
        RECT 3444.405 2631.390 3444.735 3195.910 ;
      LAYER met4 ;
        RECT 3445.135 3164.670 3588.000 3196.310 ;
        RECT 3445.135 3164.030 3445.835 3164.670 ;
        RECT 3445.135 2634.000 3445.835 3163.000 ;
        RECT 3445.135 2632.330 3445.835 2633.035 ;
      LAYER met4 ;
        RECT 3446.235 2632.730 3450.685 3164.270 ;
      LAYER met4 ;
        RECT 3451.085 3164.030 3451.685 3164.670 ;
        RECT 3451.085 2634.000 3451.685 3159.000 ;
        RECT 3451.085 2632.330 3451.685 2633.035 ;
      LAYER met4 ;
        RECT 3452.085 2632.730 3456.535 3164.270 ;
      LAYER met4 ;
        RECT 3456.935 3164.030 3457.635 3164.670 ;
        RECT 3456.935 3158.000 3458.035 3163.000 ;
      LAYER met4 ;
        RECT 3458.035 3158.000 3483.000 3164.270 ;
      LAYER met4 ;
        RECT 3483.400 3164.030 3563.385 3164.670 ;
      LAYER met4 ;
        RECT 3563.785 3163.000 3588.000 3164.270 ;
      LAYER met4 ;
        RECT 3483.000 3158.000 3485.035 3163.000 ;
        RECT 3456.935 3155.000 3485.035 3158.000 ;
        RECT 3456.935 3153.000 3458.035 3155.000 ;
      LAYER met4 ;
        RECT 3458.035 3153.000 3483.000 3155.000 ;
      LAYER met4 ;
        RECT 3483.000 3153.000 3485.035 3155.000 ;
        RECT 3456.935 3135.000 3485.035 3153.000 ;
        RECT 3456.935 3133.000 3458.035 3135.000 ;
      LAYER met4 ;
        RECT 3458.035 3133.000 3483.000 3135.000 ;
      LAYER met4 ;
        RECT 3483.000 3133.000 3485.035 3135.000 ;
        RECT 3456.935 3115.000 3485.035 3133.000 ;
        RECT 3456.935 3113.000 3458.035 3115.000 ;
      LAYER met4 ;
        RECT 3458.035 3113.000 3483.000 3115.000 ;
      LAYER met4 ;
        RECT 3483.000 3113.000 3485.035 3115.000 ;
        RECT 3456.935 3095.000 3485.035 3113.000 ;
        RECT 3456.935 3093.000 3458.035 3095.000 ;
      LAYER met4 ;
        RECT 3458.035 3093.000 3483.000 3095.000 ;
      LAYER met4 ;
        RECT 3483.000 3093.000 3485.035 3095.000 ;
        RECT 3456.935 3075.000 3485.035 3093.000 ;
        RECT 3456.935 3073.000 3458.035 3075.000 ;
      LAYER met4 ;
        RECT 3458.035 3073.000 3483.000 3075.000 ;
      LAYER met4 ;
        RECT 3483.000 3073.000 3485.035 3075.000 ;
        RECT 3456.935 3055.000 3485.035 3073.000 ;
        RECT 3456.935 3053.000 3458.035 3055.000 ;
      LAYER met4 ;
        RECT 3458.035 3053.000 3483.000 3055.000 ;
      LAYER met4 ;
        RECT 3483.000 3053.000 3485.035 3055.000 ;
        RECT 3456.935 3035.000 3485.035 3053.000 ;
        RECT 3456.935 3033.000 3458.035 3035.000 ;
      LAYER met4 ;
        RECT 3458.035 3033.000 3483.000 3035.000 ;
      LAYER met4 ;
        RECT 3483.000 3033.000 3485.035 3035.000 ;
        RECT 3456.935 3015.000 3485.035 3033.000 ;
        RECT 3456.935 3013.000 3458.035 3015.000 ;
      LAYER met4 ;
        RECT 3458.035 3013.000 3483.000 3015.000 ;
      LAYER met4 ;
        RECT 3483.000 3013.000 3485.035 3015.000 ;
        RECT 3456.935 2995.000 3485.035 3013.000 ;
        RECT 3456.935 2993.000 3458.035 2995.000 ;
      LAYER met4 ;
        RECT 3458.035 2993.000 3483.000 2995.000 ;
      LAYER met4 ;
        RECT 3483.000 2993.000 3485.035 2995.000 ;
        RECT 3456.935 2975.000 3485.035 2993.000 ;
        RECT 3456.935 2973.000 3458.035 2975.000 ;
      LAYER met4 ;
        RECT 3458.035 2973.000 3483.000 2975.000 ;
      LAYER met4 ;
        RECT 3483.000 2973.000 3485.035 2975.000 ;
        RECT 3456.935 2955.000 3485.035 2973.000 ;
        RECT 3456.935 2953.000 3458.035 2955.000 ;
      LAYER met4 ;
        RECT 3458.035 2953.000 3483.000 2955.000 ;
      LAYER met4 ;
        RECT 3483.000 2953.000 3485.035 2955.000 ;
        RECT 3456.935 2935.000 3485.035 2953.000 ;
        RECT 3456.935 2933.000 3458.035 2935.000 ;
      LAYER met4 ;
        RECT 3458.035 2933.000 3483.000 2935.000 ;
      LAYER met4 ;
        RECT 3483.000 2933.000 3485.035 2935.000 ;
        RECT 3456.935 2915.000 3485.035 2933.000 ;
        RECT 3456.935 2913.000 3458.035 2915.000 ;
      LAYER met4 ;
        RECT 3458.035 2913.000 3483.000 2915.000 ;
      LAYER met4 ;
        RECT 3483.000 2913.000 3485.035 2915.000 ;
        RECT 3456.935 2895.000 3485.035 2913.000 ;
        RECT 3456.935 2893.000 3458.035 2895.000 ;
      LAYER met4 ;
        RECT 3458.035 2893.000 3483.000 2895.000 ;
      LAYER met4 ;
        RECT 3483.000 2893.000 3485.035 2895.000 ;
        RECT 3456.935 2875.000 3485.035 2893.000 ;
        RECT 3456.935 2873.000 3458.035 2875.000 ;
      LAYER met4 ;
        RECT 3458.035 2873.000 3483.000 2875.000 ;
      LAYER met4 ;
        RECT 3483.000 2873.000 3485.035 2875.000 ;
        RECT 3456.935 2855.000 3485.035 2873.000 ;
        RECT 3456.935 2853.000 3458.035 2855.000 ;
      LAYER met4 ;
        RECT 3458.035 2853.000 3483.000 2855.000 ;
      LAYER met4 ;
        RECT 3483.000 2853.000 3485.035 2855.000 ;
        RECT 3456.935 2835.000 3485.035 2853.000 ;
        RECT 3456.935 2833.000 3458.035 2835.000 ;
      LAYER met4 ;
        RECT 3458.035 2833.000 3483.000 2835.000 ;
      LAYER met4 ;
        RECT 3483.000 2833.000 3485.035 2835.000 ;
        RECT 3456.935 2815.000 3485.035 2833.000 ;
        RECT 3456.935 2813.000 3458.035 2815.000 ;
      LAYER met4 ;
        RECT 3458.035 2813.000 3483.000 2815.000 ;
      LAYER met4 ;
        RECT 3483.000 2813.000 3485.035 2815.000 ;
        RECT 3456.935 2795.000 3485.035 2813.000 ;
        RECT 3456.935 2793.000 3458.035 2795.000 ;
      LAYER met4 ;
        RECT 3458.035 2793.000 3483.000 2795.000 ;
      LAYER met4 ;
        RECT 3483.000 2793.000 3485.035 2795.000 ;
        RECT 3456.935 2775.000 3485.035 2793.000 ;
        RECT 3456.935 2773.000 3458.035 2775.000 ;
      LAYER met4 ;
        RECT 3458.035 2773.000 3483.000 2775.000 ;
      LAYER met4 ;
        RECT 3483.000 2773.000 3485.035 2775.000 ;
        RECT 3456.935 2755.000 3485.035 2773.000 ;
        RECT 3456.935 2753.000 3458.035 2755.000 ;
      LAYER met4 ;
        RECT 3458.035 2753.000 3483.000 2755.000 ;
      LAYER met4 ;
        RECT 3483.000 2753.000 3485.035 2755.000 ;
        RECT 3456.935 2735.000 3485.035 2753.000 ;
        RECT 3456.935 2733.000 3458.035 2735.000 ;
      LAYER met4 ;
        RECT 3458.035 2733.000 3483.000 2735.000 ;
      LAYER met4 ;
        RECT 3483.000 2733.000 3485.035 2735.000 ;
        RECT 3456.935 2715.000 3485.035 2733.000 ;
        RECT 3456.935 2713.000 3458.035 2715.000 ;
      LAYER met4 ;
        RECT 3458.035 2713.000 3483.000 2715.000 ;
      LAYER met4 ;
        RECT 3483.000 2713.000 3485.035 2715.000 ;
        RECT 3456.935 2695.000 3485.035 2713.000 ;
        RECT 3456.935 2693.000 3458.035 2695.000 ;
      LAYER met4 ;
        RECT 3458.035 2693.000 3483.000 2695.000 ;
      LAYER met4 ;
        RECT 3483.000 2693.000 3485.035 2695.000 ;
        RECT 3456.935 2675.000 3485.035 2693.000 ;
        RECT 3456.935 2673.000 3458.035 2675.000 ;
      LAYER met4 ;
        RECT 3458.035 2673.000 3483.000 2675.000 ;
      LAYER met4 ;
        RECT 3483.000 2673.000 3485.035 2675.000 ;
        RECT 3456.935 2655.000 3485.035 2673.000 ;
        RECT 3456.935 2653.000 3458.035 2655.000 ;
      LAYER met4 ;
        RECT 3458.035 2653.000 3483.000 2655.000 ;
      LAYER met4 ;
        RECT 3483.000 2653.000 3485.035 2655.000 ;
        RECT 3456.935 2635.000 3485.035 2653.000 ;
        RECT 3456.935 2634.000 3458.035 2635.000 ;
        RECT 3456.935 2632.330 3457.635 2633.035 ;
      LAYER met4 ;
        RECT 3458.035 2632.730 3483.000 2635.000 ;
      LAYER met4 ;
        RECT 3483.000 2634.000 3485.035 2635.000 ;
        RECT 3562.035 2634.000 3588.000 3163.000 ;
        RECT 3483.400 2632.330 3563.385 2633.035 ;
      LAYER met4 ;
        RECT 3563.785 2632.730 3588.000 2634.000 ;
      LAYER met4 ;
        RECT 3445.135 2630.990 3588.000 2632.330 ;
        RECT 3444.505 2597.160 3588.000 2630.990 ;
        RECT 3439.745 2595.640 3588.000 2597.160 ;
        RECT 3439.745 2581.455 3440.725 2595.640 ;
        RECT 3436.465 2579.935 3440.725 2581.455 ;
        RECT 3388.535 1978.310 3435.965 2021.990 ;
      LAYER met4 ;
        RECT 3369.335 1932.055 3369.665 1932.385 ;
        RECT 3382.230 1865.490 3382.530 1956.550 ;
      LAYER met4 ;
        RECT 3388.535 1946.670 3435.335 1978.310 ;
        RECT 3388.535 1946.030 3389.635 1946.670 ;
      LAYER met4 ;
        RECT 3381.790 1864.310 3382.970 1865.490 ;
        RECT 3380.870 1860.910 3382.050 1862.090 ;
        RECT 223.855 1834.815 224.185 1835.145 ;
        RECT 223.870 1765.785 224.170 1834.815 ;
        RECT 3381.310 1786.850 3381.610 1860.910 ;
        RECT 3381.310 1786.550 3382.530 1786.850 ;
        RECT 223.855 1765.455 224.185 1765.785 ;
        RECT 3382.230 1763.050 3382.530 1786.550 ;
        RECT 3382.230 1762.750 3385.290 1763.050 ;
        RECT 3384.990 1671.250 3385.290 1762.750 ;
        RECT 3384.070 1670.950 3385.290 1671.250 ;
        RECT 3384.070 1579.450 3384.370 1670.950 ;
        RECT 3383.150 1579.150 3384.370 1579.450 ;
        RECT 3383.150 1569.250 3383.450 1579.150 ;
        RECT 3382.230 1568.950 3383.450 1569.250 ;
        RECT 3382.230 1531.850 3382.530 1568.950 ;
        RECT 3380.390 1531.550 3382.530 1531.850 ;
        RECT 3380.390 1436.650 3380.690 1531.550 ;
        RECT 3380.390 1436.350 3383.450 1436.650 ;
      LAYER met4 ;
        RECT 198.365 1419.330 199.465 1419.970 ;
        RECT 152.665 1387.690 199.465 1419.330 ;
        RECT 152.035 1344.010 199.465 1387.690 ;
      LAYER met4 ;
        RECT 3383.150 1351.650 3383.450 1436.350 ;
      LAYER met4 ;
        RECT 147.275 784.545 151.535 786.065 ;
        RECT 147.275 770.360 148.255 784.545 ;
        RECT 0.000 768.840 148.255 770.360 ;
        RECT 0.000 735.010 143.495 768.840 ;
        RECT 0.000 733.670 142.865 735.010 ;
      LAYER met4 ;
        RECT 0.000 732.000 24.215 733.270 ;
      LAYER met4 ;
        RECT 24.615 732.965 104.600 733.670 ;
        RECT 0.000 204.000 25.965 732.000 ;
        RECT 102.965 728.000 105.000 732.000 ;
      LAYER met4 ;
        RECT 105.000 728.000 129.965 733.270 ;
      LAYER met4 ;
        RECT 130.365 732.965 131.065 733.670 ;
        RECT 129.965 728.000 131.065 732.000 ;
        RECT 102.965 725.000 131.065 728.000 ;
        RECT 102.965 723.000 105.000 725.000 ;
      LAYER met4 ;
        RECT 105.000 723.000 129.965 725.000 ;
      LAYER met4 ;
        RECT 129.965 723.000 131.065 725.000 ;
        RECT 102.965 705.000 131.065 723.000 ;
        RECT 102.965 703.000 105.000 705.000 ;
      LAYER met4 ;
        RECT 105.000 703.000 129.965 705.000 ;
      LAYER met4 ;
        RECT 129.965 703.000 131.065 705.000 ;
        RECT 102.965 685.000 131.065 703.000 ;
        RECT 102.965 683.000 105.000 685.000 ;
      LAYER met4 ;
        RECT 105.000 683.000 129.965 685.000 ;
      LAYER met4 ;
        RECT 129.965 683.000 131.065 685.000 ;
        RECT 102.965 665.000 131.065 683.000 ;
        RECT 102.965 663.000 105.000 665.000 ;
      LAYER met4 ;
        RECT 105.000 663.000 129.965 665.000 ;
      LAYER met4 ;
        RECT 129.965 663.000 131.065 665.000 ;
        RECT 102.965 645.000 131.065 663.000 ;
        RECT 102.965 643.000 105.000 645.000 ;
      LAYER met4 ;
        RECT 105.000 643.000 129.965 645.000 ;
      LAYER met4 ;
        RECT 129.965 643.000 131.065 645.000 ;
        RECT 102.965 625.000 131.065 643.000 ;
        RECT 102.965 623.000 105.000 625.000 ;
      LAYER met4 ;
        RECT 105.000 623.000 129.965 625.000 ;
      LAYER met4 ;
        RECT 129.965 623.000 131.065 625.000 ;
        RECT 102.965 605.000 131.065 623.000 ;
        RECT 102.965 603.000 105.000 605.000 ;
      LAYER met4 ;
        RECT 105.000 603.000 129.965 605.000 ;
      LAYER met4 ;
        RECT 129.965 603.000 131.065 605.000 ;
        RECT 102.965 585.000 131.065 603.000 ;
        RECT 102.965 583.000 105.000 585.000 ;
      LAYER met4 ;
        RECT 105.000 583.000 129.965 585.000 ;
      LAYER met4 ;
        RECT 129.965 583.000 131.065 585.000 ;
        RECT 102.965 565.000 131.065 583.000 ;
        RECT 102.965 563.000 105.000 565.000 ;
      LAYER met4 ;
        RECT 105.000 563.000 129.965 565.000 ;
      LAYER met4 ;
        RECT 129.965 563.000 131.065 565.000 ;
        RECT 102.965 545.000 131.065 563.000 ;
        RECT 102.965 543.000 105.000 545.000 ;
      LAYER met4 ;
        RECT 105.000 543.000 129.965 545.000 ;
      LAYER met4 ;
        RECT 129.965 543.000 131.065 545.000 ;
        RECT 102.965 525.000 131.065 543.000 ;
        RECT 102.965 523.000 105.000 525.000 ;
      LAYER met4 ;
        RECT 105.000 523.000 129.965 525.000 ;
      LAYER met4 ;
        RECT 129.965 523.000 131.065 525.000 ;
        RECT 102.965 505.000 131.065 523.000 ;
        RECT 102.965 503.000 105.000 505.000 ;
      LAYER met4 ;
        RECT 105.000 503.000 129.965 505.000 ;
      LAYER met4 ;
        RECT 129.965 503.000 131.065 505.000 ;
        RECT 102.965 485.000 131.065 503.000 ;
        RECT 102.965 483.000 105.000 485.000 ;
      LAYER met4 ;
        RECT 105.000 483.000 129.965 485.000 ;
      LAYER met4 ;
        RECT 129.965 483.000 131.065 485.000 ;
        RECT 102.965 465.000 131.065 483.000 ;
        RECT 102.965 463.000 105.000 465.000 ;
      LAYER met4 ;
        RECT 105.000 463.000 129.965 465.000 ;
      LAYER met4 ;
        RECT 129.965 463.000 131.065 465.000 ;
        RECT 102.965 445.000 131.065 463.000 ;
        RECT 102.965 443.000 105.000 445.000 ;
      LAYER met4 ;
        RECT 105.000 443.000 129.965 445.000 ;
      LAYER met4 ;
        RECT 129.965 443.000 131.065 445.000 ;
        RECT 102.965 425.000 131.065 443.000 ;
        RECT 102.965 423.000 105.000 425.000 ;
      LAYER met4 ;
        RECT 105.000 423.000 129.965 425.000 ;
      LAYER met4 ;
        RECT 129.965 423.000 131.065 425.000 ;
        RECT 102.965 405.000 131.065 423.000 ;
        RECT 102.965 403.000 105.000 405.000 ;
      LAYER met4 ;
        RECT 105.000 403.000 129.965 405.000 ;
      LAYER met4 ;
        RECT 129.965 403.000 131.065 405.000 ;
        RECT 102.965 385.000 131.065 403.000 ;
        RECT 102.965 383.000 105.000 385.000 ;
      LAYER met4 ;
        RECT 105.000 383.000 129.965 385.000 ;
      LAYER met4 ;
        RECT 129.965 383.000 131.065 385.000 ;
        RECT 102.965 365.000 131.065 383.000 ;
        RECT 102.965 363.000 105.000 365.000 ;
      LAYER met4 ;
        RECT 105.000 363.000 129.965 365.000 ;
      LAYER met4 ;
        RECT 129.965 363.000 131.065 365.000 ;
        RECT 102.965 345.000 131.065 363.000 ;
        RECT 102.965 343.000 105.000 345.000 ;
      LAYER met4 ;
        RECT 105.000 343.000 129.965 345.000 ;
      LAYER met4 ;
        RECT 129.965 343.000 131.065 345.000 ;
        RECT 102.965 325.000 131.065 343.000 ;
        RECT 102.965 323.000 105.000 325.000 ;
      LAYER met4 ;
        RECT 105.000 323.000 129.965 325.000 ;
      LAYER met4 ;
        RECT 129.965 323.000 131.065 325.000 ;
        RECT 102.965 305.000 131.065 323.000 ;
        RECT 102.965 303.000 105.000 305.000 ;
      LAYER met4 ;
        RECT 105.000 303.000 129.965 305.000 ;
      LAYER met4 ;
        RECT 129.965 303.000 131.065 305.000 ;
        RECT 102.965 285.000 131.065 303.000 ;
        RECT 102.965 283.000 105.000 285.000 ;
      LAYER met4 ;
        RECT 105.000 283.000 129.965 285.000 ;
      LAYER met4 ;
        RECT 129.965 283.000 131.065 285.000 ;
        RECT 102.965 265.000 131.065 283.000 ;
        RECT 102.965 263.000 105.000 265.000 ;
      LAYER met4 ;
        RECT 105.000 263.000 129.965 265.000 ;
      LAYER met4 ;
        RECT 129.965 263.000 131.065 265.000 ;
        RECT 102.965 245.000 131.065 263.000 ;
        RECT 102.965 243.000 105.000 245.000 ;
      LAYER met4 ;
        RECT 105.000 243.000 129.965 245.000 ;
      LAYER met4 ;
        RECT 129.965 243.000 131.065 245.000 ;
        RECT 102.965 225.000 131.065 243.000 ;
        RECT 102.965 223.000 105.000 225.000 ;
      LAYER met4 ;
        RECT 105.000 223.000 129.965 225.000 ;
      LAYER met4 ;
        RECT 129.965 223.000 131.065 225.000 ;
        RECT 102.965 205.000 131.065 223.000 ;
        RECT 102.965 204.000 105.000 205.000 ;
      LAYER met4 ;
        RECT 0.000 202.730 24.215 204.000 ;
      LAYER met4 ;
        RECT 24.615 202.330 104.600 202.745 ;
        RECT 0.000 201.745 104.600 202.330 ;
      LAYER met4 ;
        RECT 105.000 202.145 129.965 205.000 ;
      LAYER met4 ;
        RECT 129.965 204.000 131.065 205.000 ;
        RECT 130.365 202.330 131.065 202.745 ;
      LAYER met4 ;
        RECT 131.465 202.730 135.915 733.270 ;
      LAYER met4 ;
        RECT 136.315 732.965 136.915 733.670 ;
        RECT 136.315 204.000 136.915 729.000 ;
        RECT 136.315 202.330 136.915 202.745 ;
      LAYER met4 ;
        RECT 137.315 202.730 141.765 733.270 ;
      LAYER met4 ;
        RECT 142.165 732.965 142.865 733.670 ;
        RECT 142.165 204.000 142.865 732.000 ;
        RECT 142.165 202.330 142.865 202.745 ;
        RECT 130.365 201.745 142.865 202.330 ;
        RECT 0.000 176.425 142.865 201.745 ;
      LAYER met4 ;
        RECT 143.265 176.825 143.595 734.610 ;
        RECT 143.895 177.090 146.875 768.440 ;
      LAYER met4 ;
        RECT 147.275 733.670 148.255 768.840 ;
      LAYER met4 ;
        RECT 147.175 732.000 148.355 733.270 ;
      LAYER met4 ;
        RECT 147.275 204.000 148.255 732.000 ;
      LAYER met4 ;
        RECT 147.175 182.445 148.355 204.000 ;
        RECT 148.655 183.125 151.635 784.145 ;
        RECT 151.935 779.090 152.265 1343.610 ;
      LAYER met4 ;
        RECT 152.665 1342.670 199.465 1344.010 ;
        RECT 152.665 1341.965 153.365 1342.670 ;
        RECT 152.665 810.330 153.365 810.970 ;
      LAYER met4 ;
        RECT 153.765 810.730 158.415 1342.270 ;
      LAYER met4 ;
        RECT 158.815 1341.965 159.415 1342.670 ;
        RECT 158.815 810.330 159.415 810.970 ;
      LAYER met4 ;
        RECT 159.815 810.730 163.265 1342.270 ;
      LAYER met4 ;
        RECT 163.665 1341.965 164.265 1342.670 ;
        RECT 163.665 810.330 164.265 810.970 ;
      LAYER met4 ;
        RECT 164.665 810.730 168.115 1342.270 ;
      LAYER met4 ;
        RECT 168.515 1341.965 169.115 1342.670 ;
        RECT 168.515 810.330 169.115 810.970 ;
      LAYER met4 ;
        RECT 169.515 810.730 174.165 1342.270 ;
      LAYER met4 ;
        RECT 174.565 1341.965 175.165 1342.670 ;
        RECT 180.615 1342.365 186.065 1342.670 ;
        RECT 174.565 810.330 175.165 810.970 ;
      LAYER met4 ;
        RECT 175.565 810.730 180.215 1342.270 ;
      LAYER met4 ;
        RECT 180.615 1341.965 181.215 1342.365 ;
        RECT 185.465 1341.965 186.065 1342.365 ;
      LAYER met4 ;
        RECT 181.615 810.970 185.065 1341.965 ;
      LAYER met4 ;
        RECT 180.615 810.570 181.215 810.970 ;
        RECT 185.465 810.570 186.065 810.970 ;
      LAYER met4 ;
        RECT 186.465 810.730 191.115 1342.270 ;
      LAYER met4 ;
        RECT 191.515 1341.965 192.115 1342.670 ;
        RECT 180.615 810.330 186.065 810.570 ;
        RECT 191.515 810.330 192.115 810.970 ;
      LAYER met4 ;
        RECT 192.515 810.730 197.965 1342.270 ;
      LAYER met4 ;
        RECT 198.365 1341.965 199.465 1342.670 ;
      LAYER met4 ;
        RECT 3382.230 1351.350 3383.450 1351.650 ;
      LAYER met4 ;
        RECT 3388.535 1415.330 3389.635 1416.035 ;
      LAYER met4 ;
        RECT 3390.035 1415.730 3395.485 1946.270 ;
      LAYER met4 ;
        RECT 3395.885 1946.030 3396.485 1946.670 ;
        RECT 3401.935 1946.430 3407.385 1946.670 ;
        RECT 3395.885 1415.330 3396.485 1416.035 ;
      LAYER met4 ;
        RECT 3396.885 1415.730 3401.535 1946.270 ;
      LAYER met4 ;
        RECT 3401.935 1946.030 3402.535 1946.430 ;
        RECT 3406.785 1946.030 3407.385 1946.430 ;
      LAYER met4 ;
        RECT 3402.935 1416.035 3406.385 1946.030 ;
      LAYER met4 ;
        RECT 3401.935 1415.635 3402.535 1416.035 ;
        RECT 3406.785 1415.635 3407.385 1416.035 ;
      LAYER met4 ;
        RECT 3407.785 1415.730 3412.435 1946.270 ;
      LAYER met4 ;
        RECT 3412.835 1946.030 3413.435 1946.670 ;
        RECT 3401.935 1415.330 3407.385 1415.635 ;
        RECT 3412.835 1415.330 3413.435 1416.035 ;
      LAYER met4 ;
        RECT 3413.835 1415.730 3418.485 1946.270 ;
      LAYER met4 ;
        RECT 3418.885 1946.030 3419.485 1946.670 ;
        RECT 3418.885 1415.330 3419.485 1416.035 ;
      LAYER met4 ;
        RECT 3419.885 1415.730 3423.335 1946.270 ;
      LAYER met4 ;
        RECT 3423.735 1946.030 3424.335 1946.670 ;
        RECT 3423.735 1415.330 3424.335 1416.035 ;
      LAYER met4 ;
        RECT 3424.735 1415.730 3428.185 1946.270 ;
      LAYER met4 ;
        RECT 3428.585 1946.030 3429.185 1946.670 ;
        RECT 3428.585 1415.330 3429.185 1416.035 ;
      LAYER met4 ;
        RECT 3429.585 1415.730 3434.235 1946.270 ;
      LAYER met4 ;
        RECT 3434.635 1946.030 3435.335 1946.670 ;
        RECT 3434.635 1415.330 3435.335 1416.035 ;
        RECT 3388.535 1413.990 3435.335 1415.330 ;
      LAYER met4 ;
        RECT 3435.735 1414.390 3436.065 1977.910 ;
        RECT 3436.365 1972.855 3439.345 2579.535 ;
      LAYER met4 ;
        RECT 3439.745 2555.670 3440.725 2579.935 ;
      LAYER met4 ;
        RECT 3439.645 2554.000 3440.825 2555.270 ;
      LAYER met4 ;
        RECT 3439.745 2025.000 3440.725 2554.000 ;
      LAYER met4 ;
        RECT 3439.645 2023.730 3440.825 2025.000 ;
      LAYER met4 ;
        RECT 3439.745 1988.160 3440.725 2023.330 ;
      LAYER met4 ;
        RECT 3441.125 1988.560 3444.105 2595.240 ;
      LAYER met4 ;
        RECT 3444.505 2587.310 3588.000 2595.640 ;
      LAYER met4 ;
        RECT 3444.405 2022.390 3444.735 2586.910 ;
      LAYER met4 ;
        RECT 3445.135 2555.670 3588.000 2587.310 ;
        RECT 3445.135 2555.030 3445.835 2555.670 ;
        RECT 3445.135 2025.000 3445.835 2554.000 ;
        RECT 3445.135 2023.330 3445.835 2024.035 ;
      LAYER met4 ;
        RECT 3446.235 2023.730 3450.685 2555.270 ;
      LAYER met4 ;
        RECT 3451.085 2555.030 3451.685 2555.670 ;
        RECT 3451.085 2025.000 3451.685 2550.000 ;
        RECT 3451.085 2023.330 3451.685 2024.035 ;
      LAYER met4 ;
        RECT 3452.085 2023.730 3456.535 2555.270 ;
      LAYER met4 ;
        RECT 3456.935 2555.030 3457.635 2555.670 ;
        RECT 3456.935 2549.000 3458.035 2554.000 ;
      LAYER met4 ;
        RECT 3458.035 2549.000 3483.000 2555.270 ;
      LAYER met4 ;
        RECT 3483.400 2555.030 3563.385 2555.670 ;
      LAYER met4 ;
        RECT 3563.785 2554.000 3588.000 2555.270 ;
      LAYER met4 ;
        RECT 3483.000 2549.000 3485.035 2554.000 ;
        RECT 3456.935 2546.000 3485.035 2549.000 ;
        RECT 3456.935 2544.000 3458.035 2546.000 ;
      LAYER met4 ;
        RECT 3458.035 2544.000 3483.000 2546.000 ;
      LAYER met4 ;
        RECT 3483.000 2544.000 3485.035 2546.000 ;
        RECT 3456.935 2526.000 3485.035 2544.000 ;
        RECT 3456.935 2524.000 3458.035 2526.000 ;
      LAYER met4 ;
        RECT 3458.035 2524.000 3483.000 2526.000 ;
      LAYER met4 ;
        RECT 3483.000 2524.000 3485.035 2526.000 ;
        RECT 3456.935 2506.000 3485.035 2524.000 ;
        RECT 3456.935 2504.000 3458.035 2506.000 ;
      LAYER met4 ;
        RECT 3458.035 2504.000 3483.000 2506.000 ;
      LAYER met4 ;
        RECT 3483.000 2504.000 3485.035 2506.000 ;
        RECT 3456.935 2486.000 3485.035 2504.000 ;
        RECT 3456.935 2484.000 3458.035 2486.000 ;
      LAYER met4 ;
        RECT 3458.035 2484.000 3483.000 2486.000 ;
      LAYER met4 ;
        RECT 3483.000 2484.000 3485.035 2486.000 ;
        RECT 3456.935 2466.000 3485.035 2484.000 ;
        RECT 3456.935 2464.000 3458.035 2466.000 ;
      LAYER met4 ;
        RECT 3458.035 2464.000 3483.000 2466.000 ;
      LAYER met4 ;
        RECT 3483.000 2464.000 3485.035 2466.000 ;
        RECT 3456.935 2446.000 3485.035 2464.000 ;
        RECT 3456.935 2444.000 3458.035 2446.000 ;
      LAYER met4 ;
        RECT 3458.035 2444.000 3483.000 2446.000 ;
      LAYER met4 ;
        RECT 3483.000 2444.000 3485.035 2446.000 ;
        RECT 3456.935 2426.000 3485.035 2444.000 ;
        RECT 3456.935 2424.000 3458.035 2426.000 ;
      LAYER met4 ;
        RECT 3458.035 2424.000 3483.000 2426.000 ;
      LAYER met4 ;
        RECT 3483.000 2424.000 3485.035 2426.000 ;
        RECT 3456.935 2406.000 3485.035 2424.000 ;
        RECT 3456.935 2404.000 3458.035 2406.000 ;
      LAYER met4 ;
        RECT 3458.035 2404.000 3483.000 2406.000 ;
      LAYER met4 ;
        RECT 3483.000 2404.000 3485.035 2406.000 ;
        RECT 3456.935 2386.000 3485.035 2404.000 ;
        RECT 3456.935 2384.000 3458.035 2386.000 ;
      LAYER met4 ;
        RECT 3458.035 2384.000 3483.000 2386.000 ;
      LAYER met4 ;
        RECT 3483.000 2384.000 3485.035 2386.000 ;
        RECT 3456.935 2366.000 3485.035 2384.000 ;
        RECT 3456.935 2364.000 3458.035 2366.000 ;
      LAYER met4 ;
        RECT 3458.035 2364.000 3483.000 2366.000 ;
      LAYER met4 ;
        RECT 3483.000 2364.000 3485.035 2366.000 ;
        RECT 3456.935 2346.000 3485.035 2364.000 ;
        RECT 3456.935 2344.000 3458.035 2346.000 ;
      LAYER met4 ;
        RECT 3458.035 2344.000 3483.000 2346.000 ;
      LAYER met4 ;
        RECT 3483.000 2344.000 3485.035 2346.000 ;
        RECT 3456.935 2326.000 3485.035 2344.000 ;
        RECT 3456.935 2324.000 3458.035 2326.000 ;
      LAYER met4 ;
        RECT 3458.035 2324.000 3483.000 2326.000 ;
      LAYER met4 ;
        RECT 3483.000 2324.000 3485.035 2326.000 ;
        RECT 3456.935 2306.000 3485.035 2324.000 ;
        RECT 3456.935 2304.000 3458.035 2306.000 ;
      LAYER met4 ;
        RECT 3458.035 2304.000 3483.000 2306.000 ;
      LAYER met4 ;
        RECT 3483.000 2304.000 3485.035 2306.000 ;
        RECT 3456.935 2286.000 3485.035 2304.000 ;
        RECT 3456.935 2284.000 3458.035 2286.000 ;
      LAYER met4 ;
        RECT 3458.035 2284.000 3483.000 2286.000 ;
      LAYER met4 ;
        RECT 3483.000 2284.000 3485.035 2286.000 ;
        RECT 3456.935 2266.000 3485.035 2284.000 ;
        RECT 3456.935 2264.000 3458.035 2266.000 ;
      LAYER met4 ;
        RECT 3458.035 2264.000 3483.000 2266.000 ;
      LAYER met4 ;
        RECT 3483.000 2264.000 3485.035 2266.000 ;
        RECT 3456.935 2246.000 3485.035 2264.000 ;
        RECT 3456.935 2244.000 3458.035 2246.000 ;
      LAYER met4 ;
        RECT 3458.035 2244.000 3483.000 2246.000 ;
      LAYER met4 ;
        RECT 3483.000 2244.000 3485.035 2246.000 ;
        RECT 3456.935 2226.000 3485.035 2244.000 ;
        RECT 3456.935 2224.000 3458.035 2226.000 ;
      LAYER met4 ;
        RECT 3458.035 2224.000 3483.000 2226.000 ;
      LAYER met4 ;
        RECT 3483.000 2224.000 3485.035 2226.000 ;
        RECT 3456.935 2206.000 3485.035 2224.000 ;
        RECT 3456.935 2204.000 3458.035 2206.000 ;
      LAYER met4 ;
        RECT 3458.035 2204.000 3483.000 2206.000 ;
      LAYER met4 ;
        RECT 3483.000 2204.000 3485.035 2206.000 ;
        RECT 3456.935 2186.000 3485.035 2204.000 ;
        RECT 3456.935 2184.000 3458.035 2186.000 ;
      LAYER met4 ;
        RECT 3458.035 2184.000 3483.000 2186.000 ;
      LAYER met4 ;
        RECT 3483.000 2184.000 3485.035 2186.000 ;
        RECT 3456.935 2166.000 3485.035 2184.000 ;
        RECT 3456.935 2164.000 3458.035 2166.000 ;
      LAYER met4 ;
        RECT 3458.035 2164.000 3483.000 2166.000 ;
      LAYER met4 ;
        RECT 3483.000 2164.000 3485.035 2166.000 ;
        RECT 3456.935 2146.000 3485.035 2164.000 ;
        RECT 3456.935 2144.000 3458.035 2146.000 ;
      LAYER met4 ;
        RECT 3458.035 2144.000 3483.000 2146.000 ;
      LAYER met4 ;
        RECT 3483.000 2144.000 3485.035 2146.000 ;
        RECT 3456.935 2126.000 3485.035 2144.000 ;
        RECT 3456.935 2124.000 3458.035 2126.000 ;
      LAYER met4 ;
        RECT 3458.035 2124.000 3483.000 2126.000 ;
      LAYER met4 ;
        RECT 3483.000 2124.000 3485.035 2126.000 ;
        RECT 3456.935 2106.000 3485.035 2124.000 ;
        RECT 3456.935 2104.000 3458.035 2106.000 ;
      LAYER met4 ;
        RECT 3458.035 2104.000 3483.000 2106.000 ;
      LAYER met4 ;
        RECT 3483.000 2104.000 3485.035 2106.000 ;
        RECT 3456.935 2086.000 3485.035 2104.000 ;
        RECT 3456.935 2084.000 3458.035 2086.000 ;
      LAYER met4 ;
        RECT 3458.035 2084.000 3483.000 2086.000 ;
      LAYER met4 ;
        RECT 3483.000 2084.000 3485.035 2086.000 ;
        RECT 3456.935 2066.000 3485.035 2084.000 ;
        RECT 3456.935 2064.000 3458.035 2066.000 ;
      LAYER met4 ;
        RECT 3458.035 2064.000 3483.000 2066.000 ;
      LAYER met4 ;
        RECT 3483.000 2064.000 3485.035 2066.000 ;
        RECT 3456.935 2046.000 3485.035 2064.000 ;
        RECT 3456.935 2044.000 3458.035 2046.000 ;
      LAYER met4 ;
        RECT 3458.035 2044.000 3483.000 2046.000 ;
      LAYER met4 ;
        RECT 3483.000 2044.000 3485.035 2046.000 ;
        RECT 3456.935 2026.000 3485.035 2044.000 ;
        RECT 3456.935 2025.000 3458.035 2026.000 ;
        RECT 3456.935 2023.330 3457.635 2024.035 ;
      LAYER met4 ;
        RECT 3458.035 2023.730 3483.000 2026.000 ;
      LAYER met4 ;
        RECT 3483.000 2025.000 3485.035 2026.000 ;
        RECT 3562.035 2025.000 3588.000 2554.000 ;
        RECT 3483.400 2023.330 3563.385 2024.035 ;
      LAYER met4 ;
        RECT 3563.785 2023.730 3588.000 2025.000 ;
      LAYER met4 ;
        RECT 3445.135 2021.990 3588.000 2023.330 ;
        RECT 3444.505 1988.160 3588.000 2021.990 ;
        RECT 3439.745 1986.640 3588.000 1988.160 ;
        RECT 3439.745 1972.455 3440.725 1986.640 ;
        RECT 3436.465 1970.935 3440.725 1972.455 ;
        RECT 3388.535 1370.310 3435.965 1413.990 ;
      LAYER met4 ;
        RECT 3382.230 1338.050 3382.530 1351.350 ;
      LAYER met4 ;
        RECT 3388.535 1338.670 3435.335 1370.310 ;
      LAYER met4 ;
        RECT 3382.230 1337.750 3383.450 1338.050 ;
      LAYER met4 ;
        RECT 3388.535 1338.030 3389.635 1338.670 ;
      LAYER met4 ;
        RECT 3383.150 1242.850 3383.450 1337.750 ;
        RECT 3383.150 1242.550 3385.290 1242.850 ;
        RECT 3384.990 1185.050 3385.290 1242.550 ;
        RECT 3384.070 1184.750 3385.290 1185.050 ;
        RECT 3384.070 1089.850 3384.370 1184.750 ;
        RECT 3383.150 1089.550 3384.370 1089.850 ;
        RECT 3383.150 1015.050 3383.450 1089.550 ;
        RECT 3382.230 1014.750 3383.450 1015.050 ;
        RECT 3382.230 899.450 3382.530 1014.750 ;
        RECT 3381.310 899.150 3382.530 899.450 ;
      LAYER met4 ;
        RECT 198.365 810.330 199.465 810.970 ;
        RECT 152.665 778.690 199.465 810.330 ;
      LAYER met4 ;
        RECT 3381.310 800.850 3381.610 899.150 ;
      LAYER met4 ;
        RECT 3388.535 806.330 3389.635 807.035 ;
      LAYER met4 ;
        RECT 3390.035 806.730 3395.485 1338.270 ;
      LAYER met4 ;
        RECT 3395.885 1338.030 3396.485 1338.670 ;
        RECT 3401.935 1338.430 3407.385 1338.670 ;
        RECT 3395.885 806.330 3396.485 807.035 ;
      LAYER met4 ;
        RECT 3396.885 806.730 3401.535 1338.270 ;
      LAYER met4 ;
        RECT 3401.935 1338.030 3402.535 1338.430 ;
        RECT 3406.785 1338.030 3407.385 1338.430 ;
      LAYER met4 ;
        RECT 3402.935 807.035 3406.385 1338.030 ;
      LAYER met4 ;
        RECT 3401.935 806.635 3402.535 807.035 ;
        RECT 3406.785 806.635 3407.385 807.035 ;
      LAYER met4 ;
        RECT 3407.785 806.730 3412.435 1338.270 ;
      LAYER met4 ;
        RECT 3412.835 1338.030 3413.435 1338.670 ;
        RECT 3401.935 806.330 3407.385 806.635 ;
        RECT 3412.835 806.330 3413.435 807.035 ;
      LAYER met4 ;
        RECT 3413.835 806.730 3418.485 1338.270 ;
      LAYER met4 ;
        RECT 3418.885 1338.030 3419.485 1338.670 ;
        RECT 3418.885 806.330 3419.485 807.035 ;
      LAYER met4 ;
        RECT 3419.885 806.730 3423.335 1338.270 ;
      LAYER met4 ;
        RECT 3423.735 1338.030 3424.335 1338.670 ;
        RECT 3423.735 806.330 3424.335 807.035 ;
      LAYER met4 ;
        RECT 3424.735 806.730 3428.185 1338.270 ;
      LAYER met4 ;
        RECT 3428.585 1338.030 3429.185 1338.670 ;
        RECT 3428.585 806.330 3429.185 807.035 ;
      LAYER met4 ;
        RECT 3429.585 806.730 3434.235 1338.270 ;
      LAYER met4 ;
        RECT 3434.635 1338.030 3435.335 1338.670 ;
        RECT 3434.635 806.330 3435.335 807.035 ;
        RECT 3388.535 804.990 3435.335 806.330 ;
      LAYER met4 ;
        RECT 3435.735 805.390 3436.065 1369.910 ;
        RECT 3436.365 1364.855 3439.345 1970.535 ;
      LAYER met4 ;
        RECT 3439.745 1946.670 3440.725 1970.935 ;
      LAYER met4 ;
        RECT 3439.645 1945.000 3440.825 1946.270 ;
      LAYER met4 ;
        RECT 3439.745 1417.000 3440.725 1945.000 ;
      LAYER met4 ;
        RECT 3439.645 1415.730 3440.825 1417.000 ;
      LAYER met4 ;
        RECT 3439.745 1380.160 3440.725 1415.330 ;
      LAYER met4 ;
        RECT 3441.125 1380.560 3444.105 1986.240 ;
      LAYER met4 ;
        RECT 3444.505 1978.310 3588.000 1986.640 ;
      LAYER met4 ;
        RECT 3444.405 1414.390 3444.735 1977.910 ;
      LAYER met4 ;
        RECT 3445.135 1946.670 3588.000 1978.310 ;
        RECT 3445.135 1946.030 3445.835 1946.670 ;
        RECT 3445.135 1417.000 3445.835 1945.000 ;
        RECT 3445.135 1415.330 3445.835 1416.035 ;
      LAYER met4 ;
        RECT 3446.235 1415.730 3450.685 1946.270 ;
      LAYER met4 ;
        RECT 3451.085 1946.030 3451.685 1946.670 ;
        RECT 3451.085 1417.000 3451.685 1942.000 ;
        RECT 3451.085 1415.330 3451.685 1416.035 ;
      LAYER met4 ;
        RECT 3452.085 1415.730 3456.535 1946.270 ;
      LAYER met4 ;
        RECT 3456.935 1946.030 3457.635 1946.670 ;
        RECT 3456.935 1941.000 3458.035 1945.000 ;
      LAYER met4 ;
        RECT 3458.035 1941.000 3483.000 1946.270 ;
      LAYER met4 ;
        RECT 3483.400 1946.030 3563.385 1946.670 ;
      LAYER met4 ;
        RECT 3563.785 1945.000 3588.000 1946.270 ;
      LAYER met4 ;
        RECT 3483.000 1941.000 3485.035 1945.000 ;
        RECT 3456.935 1938.000 3485.035 1941.000 ;
        RECT 3456.935 1936.000 3458.035 1938.000 ;
      LAYER met4 ;
        RECT 3458.035 1936.000 3483.000 1938.000 ;
      LAYER met4 ;
        RECT 3483.000 1936.000 3485.035 1938.000 ;
        RECT 3456.935 1918.000 3485.035 1936.000 ;
        RECT 3456.935 1916.000 3458.035 1918.000 ;
      LAYER met4 ;
        RECT 3458.035 1916.000 3483.000 1918.000 ;
      LAYER met4 ;
        RECT 3483.000 1916.000 3485.035 1918.000 ;
        RECT 3456.935 1898.000 3485.035 1916.000 ;
        RECT 3456.935 1896.000 3458.035 1898.000 ;
      LAYER met4 ;
        RECT 3458.035 1896.000 3483.000 1898.000 ;
      LAYER met4 ;
        RECT 3483.000 1896.000 3485.035 1898.000 ;
        RECT 3456.935 1878.000 3485.035 1896.000 ;
        RECT 3456.935 1876.000 3458.035 1878.000 ;
      LAYER met4 ;
        RECT 3458.035 1876.000 3483.000 1878.000 ;
      LAYER met4 ;
        RECT 3483.000 1876.000 3485.035 1878.000 ;
        RECT 3456.935 1858.000 3485.035 1876.000 ;
        RECT 3456.935 1856.000 3458.035 1858.000 ;
      LAYER met4 ;
        RECT 3458.035 1856.000 3483.000 1858.000 ;
      LAYER met4 ;
        RECT 3483.000 1856.000 3485.035 1858.000 ;
        RECT 3456.935 1838.000 3485.035 1856.000 ;
        RECT 3456.935 1836.000 3458.035 1838.000 ;
      LAYER met4 ;
        RECT 3458.035 1836.000 3483.000 1838.000 ;
      LAYER met4 ;
        RECT 3483.000 1836.000 3485.035 1838.000 ;
        RECT 3456.935 1818.000 3485.035 1836.000 ;
        RECT 3456.935 1816.000 3458.035 1818.000 ;
      LAYER met4 ;
        RECT 3458.035 1816.000 3483.000 1818.000 ;
      LAYER met4 ;
        RECT 3483.000 1816.000 3485.035 1818.000 ;
        RECT 3456.935 1798.000 3485.035 1816.000 ;
        RECT 3456.935 1796.000 3458.035 1798.000 ;
      LAYER met4 ;
        RECT 3458.035 1796.000 3483.000 1798.000 ;
      LAYER met4 ;
        RECT 3483.000 1796.000 3485.035 1798.000 ;
        RECT 3456.935 1778.000 3485.035 1796.000 ;
        RECT 3456.935 1776.000 3458.035 1778.000 ;
      LAYER met4 ;
        RECT 3458.035 1776.000 3483.000 1778.000 ;
      LAYER met4 ;
        RECT 3483.000 1776.000 3485.035 1778.000 ;
        RECT 3456.935 1758.000 3485.035 1776.000 ;
        RECT 3456.935 1756.000 3458.035 1758.000 ;
      LAYER met4 ;
        RECT 3458.035 1756.000 3483.000 1758.000 ;
      LAYER met4 ;
        RECT 3483.000 1756.000 3485.035 1758.000 ;
        RECT 3456.935 1738.000 3485.035 1756.000 ;
        RECT 3456.935 1736.000 3458.035 1738.000 ;
      LAYER met4 ;
        RECT 3458.035 1736.000 3483.000 1738.000 ;
      LAYER met4 ;
        RECT 3483.000 1736.000 3485.035 1738.000 ;
        RECT 3456.935 1718.000 3485.035 1736.000 ;
        RECT 3456.935 1716.000 3458.035 1718.000 ;
      LAYER met4 ;
        RECT 3458.035 1716.000 3483.000 1718.000 ;
      LAYER met4 ;
        RECT 3483.000 1716.000 3485.035 1718.000 ;
        RECT 3456.935 1698.000 3485.035 1716.000 ;
        RECT 3456.935 1696.000 3458.035 1698.000 ;
      LAYER met4 ;
        RECT 3458.035 1696.000 3483.000 1698.000 ;
      LAYER met4 ;
        RECT 3483.000 1696.000 3485.035 1698.000 ;
        RECT 3456.935 1678.000 3485.035 1696.000 ;
        RECT 3456.935 1676.000 3458.035 1678.000 ;
      LAYER met4 ;
        RECT 3458.035 1676.000 3483.000 1678.000 ;
      LAYER met4 ;
        RECT 3483.000 1676.000 3485.035 1678.000 ;
        RECT 3456.935 1658.000 3485.035 1676.000 ;
        RECT 3456.935 1656.000 3458.035 1658.000 ;
      LAYER met4 ;
        RECT 3458.035 1656.000 3483.000 1658.000 ;
      LAYER met4 ;
        RECT 3483.000 1656.000 3485.035 1658.000 ;
        RECT 3456.935 1638.000 3485.035 1656.000 ;
        RECT 3456.935 1636.000 3458.035 1638.000 ;
      LAYER met4 ;
        RECT 3458.035 1636.000 3483.000 1638.000 ;
      LAYER met4 ;
        RECT 3483.000 1636.000 3485.035 1638.000 ;
        RECT 3456.935 1618.000 3485.035 1636.000 ;
        RECT 3456.935 1616.000 3458.035 1618.000 ;
      LAYER met4 ;
        RECT 3458.035 1616.000 3483.000 1618.000 ;
      LAYER met4 ;
        RECT 3483.000 1616.000 3485.035 1618.000 ;
        RECT 3456.935 1598.000 3485.035 1616.000 ;
        RECT 3456.935 1596.000 3458.035 1598.000 ;
      LAYER met4 ;
        RECT 3458.035 1596.000 3483.000 1598.000 ;
      LAYER met4 ;
        RECT 3483.000 1596.000 3485.035 1598.000 ;
        RECT 3456.935 1578.000 3485.035 1596.000 ;
        RECT 3456.935 1576.000 3458.035 1578.000 ;
      LAYER met4 ;
        RECT 3458.035 1576.000 3483.000 1578.000 ;
      LAYER met4 ;
        RECT 3483.000 1576.000 3485.035 1578.000 ;
        RECT 3456.935 1558.000 3485.035 1576.000 ;
        RECT 3456.935 1556.000 3458.035 1558.000 ;
      LAYER met4 ;
        RECT 3458.035 1556.000 3483.000 1558.000 ;
      LAYER met4 ;
        RECT 3483.000 1556.000 3485.035 1558.000 ;
        RECT 3456.935 1538.000 3485.035 1556.000 ;
        RECT 3456.935 1536.000 3458.035 1538.000 ;
      LAYER met4 ;
        RECT 3458.035 1536.000 3483.000 1538.000 ;
      LAYER met4 ;
        RECT 3483.000 1536.000 3485.035 1538.000 ;
        RECT 3456.935 1518.000 3485.035 1536.000 ;
        RECT 3456.935 1516.000 3458.035 1518.000 ;
      LAYER met4 ;
        RECT 3458.035 1516.000 3483.000 1518.000 ;
      LAYER met4 ;
        RECT 3483.000 1516.000 3485.035 1518.000 ;
        RECT 3456.935 1498.000 3485.035 1516.000 ;
        RECT 3456.935 1496.000 3458.035 1498.000 ;
      LAYER met4 ;
        RECT 3458.035 1496.000 3483.000 1498.000 ;
      LAYER met4 ;
        RECT 3483.000 1496.000 3485.035 1498.000 ;
        RECT 3456.935 1478.000 3485.035 1496.000 ;
        RECT 3456.935 1476.000 3458.035 1478.000 ;
      LAYER met4 ;
        RECT 3458.035 1476.000 3483.000 1478.000 ;
      LAYER met4 ;
        RECT 3483.000 1476.000 3485.035 1478.000 ;
        RECT 3456.935 1458.000 3485.035 1476.000 ;
        RECT 3456.935 1456.000 3458.035 1458.000 ;
      LAYER met4 ;
        RECT 3458.035 1456.000 3483.000 1458.000 ;
      LAYER met4 ;
        RECT 3483.000 1456.000 3485.035 1458.000 ;
        RECT 3456.935 1438.000 3485.035 1456.000 ;
        RECT 3456.935 1436.000 3458.035 1438.000 ;
      LAYER met4 ;
        RECT 3458.035 1436.000 3483.000 1438.000 ;
      LAYER met4 ;
        RECT 3483.000 1436.000 3485.035 1438.000 ;
        RECT 3456.935 1418.000 3485.035 1436.000 ;
        RECT 3456.935 1417.000 3458.035 1418.000 ;
        RECT 3456.935 1415.330 3457.635 1416.035 ;
      LAYER met4 ;
        RECT 3458.035 1415.730 3483.000 1418.000 ;
      LAYER met4 ;
        RECT 3483.000 1417.000 3485.035 1418.000 ;
        RECT 3562.035 1417.000 3588.000 1945.000 ;
        RECT 3483.400 1415.330 3563.385 1416.035 ;
      LAYER met4 ;
        RECT 3563.785 1415.730 3588.000 1417.000 ;
      LAYER met4 ;
        RECT 3445.135 1413.990 3588.000 1415.330 ;
        RECT 3444.505 1380.160 3588.000 1413.990 ;
        RECT 3439.745 1378.640 3588.000 1380.160 ;
        RECT 3439.745 1364.455 3440.725 1378.640 ;
        RECT 3436.465 1362.935 3440.725 1364.455 ;
      LAYER met4 ;
        RECT 3381.310 800.550 3383.450 800.850 ;
      LAYER met4 ;
        RECT 152.035 735.010 199.465 778.690 ;
        RECT 148.755 182.045 151.535 182.725 ;
        RECT 147.275 180.025 151.535 182.045 ;
      LAYER met4 ;
        RECT 151.935 180.425 152.265 734.610 ;
      LAYER met4 ;
        RECT 152.665 733.670 199.465 735.010 ;
        RECT 152.665 732.965 153.365 733.670 ;
        RECT 152.665 202.330 153.365 202.745 ;
      LAYER met4 ;
        RECT 153.765 202.730 158.415 733.270 ;
      LAYER met4 ;
        RECT 158.815 732.965 159.415 733.670 ;
        RECT 158.815 202.330 159.415 202.745 ;
      LAYER met4 ;
        RECT 159.815 202.730 163.265 733.270 ;
      LAYER met4 ;
        RECT 163.665 732.965 164.265 733.670 ;
        RECT 163.665 202.330 164.265 202.745 ;
      LAYER met4 ;
        RECT 164.665 202.730 168.115 733.270 ;
      LAYER met4 ;
        RECT 168.515 732.965 169.115 733.670 ;
        RECT 168.515 202.330 169.115 202.745 ;
      LAYER met4 ;
        RECT 169.515 202.730 174.165 733.270 ;
      LAYER met4 ;
        RECT 174.565 732.965 175.165 733.670 ;
        RECT 180.615 733.365 186.065 733.670 ;
        RECT 174.565 202.330 175.165 202.745 ;
      LAYER met4 ;
        RECT 175.565 202.730 180.215 733.270 ;
      LAYER met4 ;
        RECT 180.615 732.965 181.215 733.365 ;
        RECT 185.465 732.965 186.065 733.365 ;
      LAYER met4 ;
        RECT 181.615 202.745 185.065 732.965 ;
      LAYER met4 ;
        RECT 180.615 202.345 181.215 202.745 ;
        RECT 185.465 202.345 186.065 202.745 ;
      LAYER met4 ;
        RECT 186.465 202.730 191.115 733.270 ;
      LAYER met4 ;
        RECT 191.515 732.965 192.115 733.670 ;
        RECT 180.615 202.330 186.065 202.345 ;
        RECT 191.515 202.330 192.115 202.745 ;
      LAYER met4 ;
        RECT 192.515 202.730 197.965 733.270 ;
      LAYER met4 ;
        RECT 198.365 732.965 199.465 733.670 ;
      LAYER met4 ;
        RECT 3383.150 607.050 3383.450 800.550 ;
      LAYER met4 ;
        RECT 3388.535 761.310 3435.965 804.990 ;
        RECT 3388.535 729.670 3435.335 761.310 ;
        RECT 3388.535 729.030 3389.635 729.670 ;
      LAYER met4 ;
        RECT 3381.310 606.750 3383.450 607.050 ;
        RECT 3381.310 510.505 3381.610 606.750 ;
        RECT 3381.295 510.175 3381.625 510.505 ;
        RECT 3384.975 510.175 3385.305 510.505 ;
        RECT 3384.990 482.625 3385.290 510.175 ;
        RECT 3384.975 482.295 3385.305 482.625 ;
        RECT 3384.055 386.415 3384.385 386.745 ;
        RECT 3384.070 386.065 3384.370 386.415 ;
        RECT 223.855 385.735 224.185 386.065 ;
        RECT 3384.055 385.735 3384.385 386.065 ;
        RECT 223.870 290.185 224.170 385.735 ;
        RECT 223.855 289.855 224.185 290.185 ;
        RECT 3383.135 289.855 3383.465 290.185 ;
        RECT 3383.150 221.505 3383.450 289.855 ;
        RECT 3383.135 221.175 3383.465 221.505 ;
      LAYER met4 ;
        RECT 198.365 202.330 200.000 202.745 ;
        RECT 152.665 198.365 200.000 202.330 ;
        RECT 1753.030 198.365 1831.035 199.465 ;
        RECT 3385.255 198.365 3389.635 200.000 ;
        RECT 152.665 192.115 197.250 198.365 ;
      LAYER met4 ;
        RECT 197.650 192.515 668.270 197.965 ;
      LAYER met4 ;
        RECT 668.670 192.115 740.330 197.965 ;
      LAYER met4 ;
        RECT 740.730 192.515 1209.000 197.965 ;
      LAYER met4 ;
        RECT 152.665 191.515 200.000 192.115 ;
        RECT 667.965 191.515 741.035 192.115 ;
        RECT 152.665 186.065 195.815 191.515 ;
      LAYER met4 ;
        RECT 196.215 186.465 668.270 191.115 ;
      LAYER met4 ;
        RECT 668.670 186.065 740.330 191.515 ;
      LAYER met4 ;
        RECT 740.730 186.465 1209.000 191.115 ;
      LAYER met4 ;
        RECT 152.665 185.465 200.000 186.065 ;
        RECT 667.965 185.465 741.035 186.065 ;
        RECT 152.665 181.215 198.130 185.465 ;
      LAYER met4 ;
        RECT 198.530 181.615 667.965 185.065 ;
      LAYER met4 ;
        RECT 668.365 181.215 740.635 185.465 ;
      LAYER met4 ;
        RECT 741.035 181.615 1209.000 185.065 ;
      LAYER met4 ;
        RECT 152.665 180.615 200.000 181.215 ;
        RECT 667.965 180.615 741.035 181.215 ;
        RECT 152.665 180.025 198.075 180.615 ;
        RECT 147.275 176.690 198.075 180.025 ;
        RECT 143.995 176.425 198.075 176.690 ;
        RECT 0.000 175.165 198.075 176.425 ;
      LAYER met4 ;
        RECT 198.475 175.565 668.270 180.215 ;
      LAYER met4 ;
        RECT 668.670 175.165 740.330 180.615 ;
      LAYER met4 ;
        RECT 740.730 175.565 1209.000 180.215 ;
      LAYER met4 ;
        RECT 0.000 174.565 200.000 175.165 ;
        RECT 667.965 174.565 741.035 175.165 ;
        RECT 0.000 169.115 198.000 174.565 ;
      LAYER met4 ;
        RECT 198.400 169.515 668.270 174.165 ;
      LAYER met4 ;
        RECT 668.670 169.115 740.330 174.565 ;
      LAYER met4 ;
        RECT 740.730 169.515 1209.000 174.165 ;
      LAYER met4 ;
        RECT 0.000 168.515 200.000 169.115 ;
        RECT 667.965 168.515 741.035 169.115 ;
        RECT 0.000 164.265 198.215 168.515 ;
      LAYER met4 ;
        RECT 198.615 164.665 668.270 168.115 ;
      LAYER met4 ;
        RECT 668.670 164.265 740.330 168.515 ;
      LAYER met4 ;
        RECT 740.730 164.665 1209.000 168.115 ;
      LAYER met4 ;
        RECT 0.000 163.665 200.000 164.265 ;
        RECT 667.965 163.665 741.035 164.265 ;
        RECT 0.000 159.415 198.265 163.665 ;
      LAYER met4 ;
        RECT 198.665 159.815 668.270 163.265 ;
      LAYER met4 ;
        RECT 668.670 159.415 740.330 163.665 ;
      LAYER met4 ;
        RECT 740.730 159.815 1209.000 163.265 ;
      LAYER met4 ;
        RECT 0.000 158.815 200.000 159.415 ;
        RECT 667.965 158.815 741.035 159.415 ;
        RECT 0.000 153.365 198.125 158.815 ;
      LAYER met4 ;
        RECT 198.525 153.765 668.270 158.415 ;
      LAYER met4 ;
        RECT 668.670 153.365 740.330 158.815 ;
      LAYER met4 ;
        RECT 740.730 153.765 1209.000 158.415 ;
      LAYER met4 ;
        RECT 0.000 152.665 200.000 153.365 ;
        RECT 667.965 152.665 741.035 153.365 ;
        RECT 0.000 152.035 180.025 152.665 ;
        RECT 0.000 148.755 178.665 152.035 ;
      LAYER met4 ;
        RECT 180.425 151.935 668.270 152.265 ;
      LAYER met4 ;
        RECT 668.670 152.035 740.330 152.665 ;
      LAYER met4 ;
        RECT 740.730 151.935 1209.000 152.265 ;
      LAYER met4 ;
        RECT 1209.000 152.035 1284.000 197.965 ;
      LAYER met4 ;
        RECT 1284.000 192.515 1753.270 197.965 ;
      LAYER met4 ;
        RECT 1753.670 192.115 1830.330 198.365 ;
      LAYER met4 ;
        RECT 1830.730 192.515 2300.270 197.965 ;
      LAYER met4 ;
        RECT 2300.670 192.115 2372.330 197.965 ;
      LAYER met4 ;
        RECT 2372.730 192.515 2842.270 197.965 ;
      LAYER met4 ;
        RECT 2842.670 192.115 2914.330 197.965 ;
      LAYER met4 ;
        RECT 2914.730 192.515 3385.270 197.965 ;
      LAYER met4 ;
        RECT 3385.670 197.250 3389.635 198.365 ;
      LAYER met4 ;
        RECT 3390.035 197.650 3395.485 729.270 ;
      LAYER met4 ;
        RECT 3395.885 729.030 3396.485 729.670 ;
        RECT 3401.935 729.430 3407.385 729.670 ;
        RECT 3395.885 197.250 3396.485 200.000 ;
        RECT 3385.670 195.815 3396.485 197.250 ;
      LAYER met4 ;
        RECT 3396.885 196.215 3401.535 729.270 ;
      LAYER met4 ;
        RECT 3401.935 729.030 3402.535 729.430 ;
        RECT 3406.785 729.030 3407.385 729.430 ;
        RECT 3401.935 198.130 3402.535 200.000 ;
      LAYER met4 ;
        RECT 3402.935 198.530 3406.385 729.030 ;
      LAYER met4 ;
        RECT 3406.785 198.130 3407.385 200.000 ;
      LAYER met4 ;
        RECT 3407.785 198.475 3412.435 729.270 ;
      LAYER met4 ;
        RECT 3412.835 729.030 3413.435 729.670 ;
        RECT 3401.935 198.075 3407.385 198.130 ;
        RECT 3412.835 198.075 3413.435 200.000 ;
      LAYER met4 ;
        RECT 3413.835 198.400 3418.485 729.270 ;
      LAYER met4 ;
        RECT 3418.885 729.030 3419.485 729.670 ;
        RECT 3401.935 198.000 3413.435 198.075 ;
        RECT 3418.885 198.215 3419.485 200.000 ;
      LAYER met4 ;
        RECT 3419.885 198.615 3423.335 729.270 ;
      LAYER met4 ;
        RECT 3423.735 729.030 3424.335 729.670 ;
        RECT 3423.735 198.265 3424.335 200.000 ;
      LAYER met4 ;
        RECT 3424.735 198.665 3428.185 729.270 ;
      LAYER met4 ;
        RECT 3428.585 729.030 3429.185 729.670 ;
        RECT 3428.585 198.265 3429.185 200.000 ;
      LAYER met4 ;
        RECT 3429.585 198.525 3434.235 729.270 ;
      LAYER met4 ;
        RECT 3434.635 729.030 3435.335 729.670 ;
        RECT 3423.735 198.215 3429.185 198.265 ;
        RECT 3418.885 198.125 3429.185 198.215 ;
        RECT 3434.635 198.125 3435.335 200.000 ;
        RECT 3418.885 198.000 3435.335 198.125 ;
        RECT 3401.935 195.815 3435.335 198.000 ;
        RECT 3385.670 192.115 3435.335 195.815 ;
        RECT 1753.030 191.515 1831.035 192.115 ;
        RECT 2299.965 191.515 2373.035 192.115 ;
        RECT 2841.965 191.515 2915.035 192.115 ;
        RECT 3385.255 191.515 3435.335 192.115 ;
      LAYER met4 ;
        RECT 1284.000 186.465 1753.270 191.115 ;
      LAYER met4 ;
        RECT 1753.670 186.065 1830.330 191.515 ;
      LAYER met4 ;
        RECT 1830.730 186.465 2300.270 191.115 ;
      LAYER met4 ;
        RECT 2300.670 186.065 2372.330 191.515 ;
      LAYER met4 ;
        RECT 2372.730 186.465 2842.270 191.115 ;
      LAYER met4 ;
        RECT 2842.670 186.065 2914.330 191.515 ;
      LAYER met4 ;
        RECT 2914.730 186.465 3385.270 191.115 ;
      LAYER met4 ;
        RECT 3385.670 186.065 3435.335 191.515 ;
        RECT 1753.030 185.465 1831.035 186.065 ;
        RECT 2299.965 185.465 2373.035 186.065 ;
        RECT 2841.965 185.465 2915.035 186.065 ;
        RECT 3385.255 185.465 3435.335 186.065 ;
      LAYER met4 ;
        RECT 1284.000 181.615 1753.030 185.065 ;
      LAYER met4 ;
        RECT 1753.430 181.215 1830.635 185.465 ;
      LAYER met4 ;
        RECT 1831.035 181.615 2299.965 185.065 ;
      LAYER met4 ;
        RECT 2300.365 181.215 2372.635 185.465 ;
      LAYER met4 ;
        RECT 2373.035 181.615 2841.965 185.065 ;
      LAYER met4 ;
        RECT 2842.365 181.215 2914.635 185.465 ;
      LAYER met4 ;
        RECT 2915.035 181.615 3385.255 185.065 ;
      LAYER met4 ;
        RECT 3385.655 181.215 3435.335 185.465 ;
        RECT 1753.030 180.615 1831.035 181.215 ;
        RECT 2299.965 180.615 2373.035 181.215 ;
        RECT 2841.965 180.615 2915.035 181.215 ;
        RECT 3385.255 180.615 3435.335 181.215 ;
      LAYER met4 ;
        RECT 1284.000 175.565 1753.270 180.215 ;
      LAYER met4 ;
        RECT 1753.670 175.165 1830.330 180.615 ;
      LAYER met4 ;
        RECT 1830.730 175.565 2300.270 180.215 ;
      LAYER met4 ;
        RECT 2300.670 175.165 2372.330 180.615 ;
      LAYER met4 ;
        RECT 2372.730 175.565 2842.270 180.215 ;
      LAYER met4 ;
        RECT 2842.670 175.165 2914.330 180.615 ;
      LAYER met4 ;
        RECT 2914.730 175.565 3385.270 180.215 ;
      LAYER met4 ;
        RECT 3385.670 180.025 3435.335 180.615 ;
      LAYER met4 ;
        RECT 3435.735 180.425 3436.065 760.910 ;
        RECT 3436.365 755.855 3439.345 1362.535 ;
      LAYER met4 ;
        RECT 3439.745 1338.670 3440.725 1362.935 ;
      LAYER met4 ;
        RECT 3439.645 1337.000 3440.825 1338.270 ;
      LAYER met4 ;
        RECT 3439.745 808.000 3440.725 1337.000 ;
      LAYER met4 ;
        RECT 3439.645 806.730 3440.825 808.000 ;
      LAYER met4 ;
        RECT 3439.745 771.160 3440.725 806.330 ;
      LAYER met4 ;
        RECT 3441.125 771.560 3444.105 1378.240 ;
      LAYER met4 ;
        RECT 3444.505 1370.310 3588.000 1378.640 ;
      LAYER met4 ;
        RECT 3444.405 805.390 3444.735 1369.910 ;
      LAYER met4 ;
        RECT 3445.135 1338.670 3588.000 1370.310 ;
        RECT 3445.135 1338.030 3445.835 1338.670 ;
        RECT 3445.135 808.000 3445.835 1337.000 ;
        RECT 3445.135 806.330 3445.835 807.035 ;
      LAYER met4 ;
        RECT 3446.235 806.730 3450.685 1338.270 ;
      LAYER met4 ;
        RECT 3451.085 1338.030 3451.685 1338.670 ;
        RECT 3451.085 808.000 3451.685 1333.000 ;
        RECT 3451.085 806.330 3451.685 807.035 ;
      LAYER met4 ;
        RECT 3452.085 806.730 3456.535 1338.270 ;
      LAYER met4 ;
        RECT 3456.935 1338.030 3457.635 1338.670 ;
        RECT 3456.935 1332.000 3458.035 1337.000 ;
      LAYER met4 ;
        RECT 3458.035 1332.000 3483.000 1338.270 ;
      LAYER met4 ;
        RECT 3483.400 1338.030 3563.385 1338.670 ;
      LAYER met4 ;
        RECT 3563.785 1337.000 3588.000 1338.270 ;
      LAYER met4 ;
        RECT 3483.000 1332.000 3485.035 1337.000 ;
        RECT 3456.935 1329.000 3485.035 1332.000 ;
        RECT 3456.935 1327.000 3458.035 1329.000 ;
      LAYER met4 ;
        RECT 3458.035 1327.000 3483.000 1329.000 ;
      LAYER met4 ;
        RECT 3483.000 1327.000 3485.035 1329.000 ;
        RECT 3456.935 1309.000 3485.035 1327.000 ;
        RECT 3456.935 1307.000 3458.035 1309.000 ;
      LAYER met4 ;
        RECT 3458.035 1307.000 3483.000 1309.000 ;
      LAYER met4 ;
        RECT 3483.000 1307.000 3485.035 1309.000 ;
        RECT 3456.935 1289.000 3485.035 1307.000 ;
        RECT 3456.935 1287.000 3458.035 1289.000 ;
      LAYER met4 ;
        RECT 3458.035 1287.000 3483.000 1289.000 ;
      LAYER met4 ;
        RECT 3483.000 1287.000 3485.035 1289.000 ;
        RECT 3456.935 1269.000 3485.035 1287.000 ;
        RECT 3456.935 1267.000 3458.035 1269.000 ;
      LAYER met4 ;
        RECT 3458.035 1267.000 3483.000 1269.000 ;
      LAYER met4 ;
        RECT 3483.000 1267.000 3485.035 1269.000 ;
        RECT 3456.935 1249.000 3485.035 1267.000 ;
        RECT 3456.935 1247.000 3458.035 1249.000 ;
      LAYER met4 ;
        RECT 3458.035 1247.000 3483.000 1249.000 ;
      LAYER met4 ;
        RECT 3483.000 1247.000 3485.035 1249.000 ;
        RECT 3456.935 1229.000 3485.035 1247.000 ;
        RECT 3456.935 1227.000 3458.035 1229.000 ;
      LAYER met4 ;
        RECT 3458.035 1227.000 3483.000 1229.000 ;
      LAYER met4 ;
        RECT 3483.000 1227.000 3485.035 1229.000 ;
        RECT 3456.935 1209.000 3485.035 1227.000 ;
        RECT 3456.935 1207.000 3458.035 1209.000 ;
      LAYER met4 ;
        RECT 3458.035 1207.000 3483.000 1209.000 ;
      LAYER met4 ;
        RECT 3483.000 1207.000 3485.035 1209.000 ;
        RECT 3456.935 1189.000 3485.035 1207.000 ;
        RECT 3456.935 1187.000 3458.035 1189.000 ;
      LAYER met4 ;
        RECT 3458.035 1187.000 3483.000 1189.000 ;
      LAYER met4 ;
        RECT 3483.000 1187.000 3485.035 1189.000 ;
        RECT 3456.935 1169.000 3485.035 1187.000 ;
        RECT 3456.935 1167.000 3458.035 1169.000 ;
      LAYER met4 ;
        RECT 3458.035 1167.000 3483.000 1169.000 ;
      LAYER met4 ;
        RECT 3483.000 1167.000 3485.035 1169.000 ;
        RECT 3456.935 1149.000 3485.035 1167.000 ;
        RECT 3456.935 1147.000 3458.035 1149.000 ;
      LAYER met4 ;
        RECT 3458.035 1147.000 3483.000 1149.000 ;
      LAYER met4 ;
        RECT 3483.000 1147.000 3485.035 1149.000 ;
        RECT 3456.935 1129.000 3485.035 1147.000 ;
        RECT 3456.935 1127.000 3458.035 1129.000 ;
      LAYER met4 ;
        RECT 3458.035 1127.000 3483.000 1129.000 ;
      LAYER met4 ;
        RECT 3483.000 1127.000 3485.035 1129.000 ;
        RECT 3456.935 1109.000 3485.035 1127.000 ;
        RECT 3456.935 1107.000 3458.035 1109.000 ;
      LAYER met4 ;
        RECT 3458.035 1107.000 3483.000 1109.000 ;
      LAYER met4 ;
        RECT 3483.000 1107.000 3485.035 1109.000 ;
        RECT 3456.935 1089.000 3485.035 1107.000 ;
        RECT 3456.935 1087.000 3458.035 1089.000 ;
      LAYER met4 ;
        RECT 3458.035 1087.000 3483.000 1089.000 ;
      LAYER met4 ;
        RECT 3483.000 1087.000 3485.035 1089.000 ;
        RECT 3456.935 1069.000 3485.035 1087.000 ;
        RECT 3456.935 1067.000 3458.035 1069.000 ;
      LAYER met4 ;
        RECT 3458.035 1067.000 3483.000 1069.000 ;
      LAYER met4 ;
        RECT 3483.000 1067.000 3485.035 1069.000 ;
        RECT 3456.935 1049.000 3485.035 1067.000 ;
        RECT 3456.935 1047.000 3458.035 1049.000 ;
      LAYER met4 ;
        RECT 3458.035 1047.000 3483.000 1049.000 ;
      LAYER met4 ;
        RECT 3483.000 1047.000 3485.035 1049.000 ;
        RECT 3456.935 1029.000 3485.035 1047.000 ;
        RECT 3456.935 1027.000 3458.035 1029.000 ;
      LAYER met4 ;
        RECT 3458.035 1027.000 3483.000 1029.000 ;
      LAYER met4 ;
        RECT 3483.000 1027.000 3485.035 1029.000 ;
        RECT 3456.935 1009.000 3485.035 1027.000 ;
        RECT 3456.935 1007.000 3458.035 1009.000 ;
      LAYER met4 ;
        RECT 3458.035 1007.000 3483.000 1009.000 ;
      LAYER met4 ;
        RECT 3483.000 1007.000 3485.035 1009.000 ;
        RECT 3456.935 989.000 3485.035 1007.000 ;
        RECT 3456.935 987.000 3458.035 989.000 ;
      LAYER met4 ;
        RECT 3458.035 987.000 3483.000 989.000 ;
      LAYER met4 ;
        RECT 3483.000 987.000 3485.035 989.000 ;
        RECT 3456.935 969.000 3485.035 987.000 ;
        RECT 3456.935 967.000 3458.035 969.000 ;
      LAYER met4 ;
        RECT 3458.035 967.000 3483.000 969.000 ;
      LAYER met4 ;
        RECT 3483.000 967.000 3485.035 969.000 ;
        RECT 3456.935 949.000 3485.035 967.000 ;
        RECT 3456.935 947.000 3458.035 949.000 ;
      LAYER met4 ;
        RECT 3458.035 947.000 3483.000 949.000 ;
      LAYER met4 ;
        RECT 3483.000 947.000 3485.035 949.000 ;
        RECT 3456.935 929.000 3485.035 947.000 ;
        RECT 3456.935 927.000 3458.035 929.000 ;
      LAYER met4 ;
        RECT 3458.035 927.000 3483.000 929.000 ;
      LAYER met4 ;
        RECT 3483.000 927.000 3485.035 929.000 ;
        RECT 3456.935 909.000 3485.035 927.000 ;
        RECT 3456.935 907.000 3458.035 909.000 ;
      LAYER met4 ;
        RECT 3458.035 907.000 3483.000 909.000 ;
      LAYER met4 ;
        RECT 3483.000 907.000 3485.035 909.000 ;
        RECT 3456.935 889.000 3485.035 907.000 ;
        RECT 3456.935 887.000 3458.035 889.000 ;
      LAYER met4 ;
        RECT 3458.035 887.000 3483.000 889.000 ;
      LAYER met4 ;
        RECT 3483.000 887.000 3485.035 889.000 ;
        RECT 3456.935 869.000 3485.035 887.000 ;
        RECT 3456.935 867.000 3458.035 869.000 ;
      LAYER met4 ;
        RECT 3458.035 867.000 3483.000 869.000 ;
      LAYER met4 ;
        RECT 3483.000 867.000 3485.035 869.000 ;
        RECT 3456.935 849.000 3485.035 867.000 ;
        RECT 3456.935 847.000 3458.035 849.000 ;
      LAYER met4 ;
        RECT 3458.035 847.000 3483.000 849.000 ;
      LAYER met4 ;
        RECT 3483.000 847.000 3485.035 849.000 ;
        RECT 3456.935 829.000 3485.035 847.000 ;
        RECT 3456.935 827.000 3458.035 829.000 ;
      LAYER met4 ;
        RECT 3458.035 827.000 3483.000 829.000 ;
      LAYER met4 ;
        RECT 3483.000 827.000 3485.035 829.000 ;
        RECT 3456.935 809.000 3485.035 827.000 ;
        RECT 3456.935 808.000 3458.035 809.000 ;
        RECT 3456.935 806.330 3457.635 807.035 ;
      LAYER met4 ;
        RECT 3458.035 806.730 3483.000 809.000 ;
      LAYER met4 ;
        RECT 3483.000 808.000 3485.035 809.000 ;
        RECT 3562.035 808.000 3588.000 1337.000 ;
        RECT 3483.400 806.330 3563.385 807.035 ;
      LAYER met4 ;
        RECT 3563.785 806.730 3588.000 808.000 ;
      LAYER met4 ;
        RECT 3445.135 804.990 3588.000 806.330 ;
        RECT 3444.505 771.160 3588.000 804.990 ;
        RECT 3439.745 769.640 3588.000 771.160 ;
        RECT 3439.745 755.455 3440.725 769.640 ;
        RECT 3436.465 753.935 3440.725 755.455 ;
        RECT 3385.670 178.665 3435.965 180.025 ;
      LAYER met4 ;
        RECT 3436.365 179.065 3439.345 753.535 ;
      LAYER met4 ;
        RECT 3439.745 729.670 3440.725 753.935 ;
      LAYER met4 ;
        RECT 3439.645 728.000 3440.825 729.270 ;
      LAYER met4 ;
        RECT 3439.745 200.000 3440.725 728.000 ;
        RECT 3385.670 178.050 3439.245 178.665 ;
      LAYER met4 ;
        RECT 3439.645 178.450 3440.825 200.000 ;
      LAYER met4 ;
        RECT 3385.670 176.690 3440.725 178.050 ;
      LAYER met4 ;
        RECT 3441.125 177.090 3444.105 769.240 ;
      LAYER met4 ;
        RECT 3444.505 761.310 3588.000 769.640 ;
      LAYER met4 ;
        RECT 3444.405 176.825 3444.735 760.910 ;
      LAYER met4 ;
        RECT 3445.135 729.670 3588.000 761.310 ;
        RECT 3445.135 729.030 3445.835 729.670 ;
        RECT 3445.135 197.975 3445.835 728.000 ;
      LAYER met4 ;
        RECT 3446.235 198.375 3450.685 729.270 ;
      LAYER met4 ;
        RECT 3451.085 729.030 3451.685 729.670 ;
        RECT 3451.085 198.120 3451.685 725.000 ;
      LAYER met4 ;
        RECT 3452.085 198.520 3456.535 729.270 ;
      LAYER met4 ;
        RECT 3456.935 729.030 3457.635 729.670 ;
        RECT 3456.935 724.000 3458.035 728.000 ;
      LAYER met4 ;
        RECT 3458.035 724.000 3483.000 729.270 ;
      LAYER met4 ;
        RECT 3483.400 729.030 3563.385 729.670 ;
      LAYER met4 ;
        RECT 3563.785 728.000 3588.000 729.270 ;
      LAYER met4 ;
        RECT 3483.000 724.000 3485.035 728.000 ;
        RECT 3456.935 721.000 3485.035 724.000 ;
        RECT 3456.935 719.000 3458.035 721.000 ;
      LAYER met4 ;
        RECT 3458.035 719.000 3483.000 721.000 ;
      LAYER met4 ;
        RECT 3483.000 719.000 3485.035 721.000 ;
        RECT 3456.935 701.000 3485.035 719.000 ;
        RECT 3456.935 699.000 3458.035 701.000 ;
      LAYER met4 ;
        RECT 3458.035 699.000 3483.000 701.000 ;
      LAYER met4 ;
        RECT 3483.000 699.000 3485.035 701.000 ;
        RECT 3456.935 681.000 3485.035 699.000 ;
        RECT 3456.935 679.000 3458.035 681.000 ;
      LAYER met4 ;
        RECT 3458.035 679.000 3483.000 681.000 ;
      LAYER met4 ;
        RECT 3483.000 679.000 3485.035 681.000 ;
        RECT 3456.935 661.000 3485.035 679.000 ;
        RECT 3456.935 659.000 3458.035 661.000 ;
      LAYER met4 ;
        RECT 3458.035 659.000 3483.000 661.000 ;
      LAYER met4 ;
        RECT 3483.000 659.000 3485.035 661.000 ;
        RECT 3456.935 641.000 3485.035 659.000 ;
        RECT 3456.935 639.000 3458.035 641.000 ;
      LAYER met4 ;
        RECT 3458.035 639.000 3483.000 641.000 ;
      LAYER met4 ;
        RECT 3483.000 639.000 3485.035 641.000 ;
        RECT 3456.935 621.000 3485.035 639.000 ;
        RECT 3456.935 619.000 3458.035 621.000 ;
      LAYER met4 ;
        RECT 3458.035 619.000 3483.000 621.000 ;
      LAYER met4 ;
        RECT 3483.000 619.000 3485.035 621.000 ;
        RECT 3456.935 601.000 3485.035 619.000 ;
        RECT 3456.935 599.000 3458.035 601.000 ;
      LAYER met4 ;
        RECT 3458.035 599.000 3483.000 601.000 ;
      LAYER met4 ;
        RECT 3483.000 599.000 3485.035 601.000 ;
        RECT 3456.935 581.000 3485.035 599.000 ;
        RECT 3456.935 579.000 3458.035 581.000 ;
      LAYER met4 ;
        RECT 3458.035 579.000 3483.000 581.000 ;
      LAYER met4 ;
        RECT 3483.000 579.000 3485.035 581.000 ;
        RECT 3456.935 561.000 3485.035 579.000 ;
        RECT 3456.935 559.000 3458.035 561.000 ;
      LAYER met4 ;
        RECT 3458.035 559.000 3483.000 561.000 ;
      LAYER met4 ;
        RECT 3483.000 559.000 3485.035 561.000 ;
        RECT 3456.935 541.000 3485.035 559.000 ;
        RECT 3456.935 539.000 3458.035 541.000 ;
      LAYER met4 ;
        RECT 3458.035 539.000 3483.000 541.000 ;
      LAYER met4 ;
        RECT 3483.000 539.000 3485.035 541.000 ;
        RECT 3456.935 521.000 3485.035 539.000 ;
        RECT 3456.935 519.000 3458.035 521.000 ;
      LAYER met4 ;
        RECT 3458.035 519.000 3483.000 521.000 ;
      LAYER met4 ;
        RECT 3483.000 519.000 3485.035 521.000 ;
        RECT 3456.935 501.000 3485.035 519.000 ;
        RECT 3456.935 499.000 3458.035 501.000 ;
      LAYER met4 ;
        RECT 3458.035 499.000 3483.000 501.000 ;
      LAYER met4 ;
        RECT 3483.000 499.000 3485.035 501.000 ;
        RECT 3456.935 481.000 3485.035 499.000 ;
        RECT 3456.935 479.000 3458.035 481.000 ;
      LAYER met4 ;
        RECT 3458.035 479.000 3483.000 481.000 ;
      LAYER met4 ;
        RECT 3483.000 479.000 3485.035 481.000 ;
        RECT 3456.935 461.000 3485.035 479.000 ;
        RECT 3456.935 459.000 3458.035 461.000 ;
      LAYER met4 ;
        RECT 3458.035 459.000 3483.000 461.000 ;
      LAYER met4 ;
        RECT 3483.000 459.000 3485.035 461.000 ;
        RECT 3456.935 441.000 3485.035 459.000 ;
        RECT 3456.935 439.000 3458.035 441.000 ;
      LAYER met4 ;
        RECT 3458.035 439.000 3483.000 441.000 ;
      LAYER met4 ;
        RECT 3483.000 439.000 3485.035 441.000 ;
        RECT 3456.935 421.000 3485.035 439.000 ;
        RECT 3456.935 419.000 3458.035 421.000 ;
      LAYER met4 ;
        RECT 3458.035 419.000 3483.000 421.000 ;
      LAYER met4 ;
        RECT 3483.000 419.000 3485.035 421.000 ;
        RECT 3456.935 401.000 3485.035 419.000 ;
        RECT 3456.935 399.000 3458.035 401.000 ;
      LAYER met4 ;
        RECT 3458.035 399.000 3483.000 401.000 ;
      LAYER met4 ;
        RECT 3483.000 399.000 3485.035 401.000 ;
        RECT 3456.935 381.000 3485.035 399.000 ;
        RECT 3456.935 379.000 3458.035 381.000 ;
      LAYER met4 ;
        RECT 3458.035 379.000 3483.000 381.000 ;
      LAYER met4 ;
        RECT 3483.000 379.000 3485.035 381.000 ;
        RECT 3456.935 361.000 3485.035 379.000 ;
        RECT 3456.935 359.000 3458.035 361.000 ;
      LAYER met4 ;
        RECT 3458.035 359.000 3483.000 361.000 ;
      LAYER met4 ;
        RECT 3483.000 359.000 3485.035 361.000 ;
        RECT 3456.935 341.000 3485.035 359.000 ;
        RECT 3456.935 339.000 3458.035 341.000 ;
      LAYER met4 ;
        RECT 3458.035 339.000 3483.000 341.000 ;
      LAYER met4 ;
        RECT 3483.000 339.000 3485.035 341.000 ;
        RECT 3456.935 321.000 3485.035 339.000 ;
        RECT 3456.935 319.000 3458.035 321.000 ;
      LAYER met4 ;
        RECT 3458.035 319.000 3483.000 321.000 ;
      LAYER met4 ;
        RECT 3483.000 319.000 3485.035 321.000 ;
        RECT 3456.935 301.000 3485.035 319.000 ;
        RECT 3456.935 299.000 3458.035 301.000 ;
      LAYER met4 ;
        RECT 3458.035 299.000 3483.000 301.000 ;
      LAYER met4 ;
        RECT 3483.000 299.000 3485.035 301.000 ;
        RECT 3456.935 281.000 3485.035 299.000 ;
        RECT 3456.935 279.000 3458.035 281.000 ;
      LAYER met4 ;
        RECT 3458.035 279.000 3483.000 281.000 ;
      LAYER met4 ;
        RECT 3483.000 279.000 3485.035 281.000 ;
        RECT 3456.935 261.000 3485.035 279.000 ;
        RECT 3456.935 259.000 3458.035 261.000 ;
      LAYER met4 ;
        RECT 3458.035 259.000 3483.000 261.000 ;
      LAYER met4 ;
        RECT 3483.000 259.000 3485.035 261.000 ;
        RECT 3456.935 241.000 3485.035 259.000 ;
        RECT 3456.935 239.000 3458.035 241.000 ;
      LAYER met4 ;
        RECT 3458.035 239.000 3483.000 241.000 ;
      LAYER met4 ;
        RECT 3483.000 239.000 3485.035 241.000 ;
        RECT 3456.935 221.000 3485.035 239.000 ;
        RECT 3456.935 219.000 3458.035 221.000 ;
      LAYER met4 ;
        RECT 3458.035 219.000 3483.000 221.000 ;
      LAYER met4 ;
        RECT 3483.000 219.000 3485.035 221.000 ;
        RECT 3456.935 201.000 3485.035 219.000 ;
        RECT 3456.935 200.000 3458.035 201.000 ;
        RECT 3456.935 198.120 3457.635 200.000 ;
        RECT 3451.085 197.975 3457.635 198.120 ;
        RECT 3445.135 196.955 3457.635 197.975 ;
      LAYER met4 ;
        RECT 3458.035 197.355 3483.000 201.000 ;
      LAYER met4 ;
        RECT 3483.000 200.000 3485.035 201.000 ;
        RECT 3562.035 200.000 3588.000 728.000 ;
        RECT 3483.400 198.165 3563.385 200.000 ;
      LAYER met4 ;
        RECT 3563.785 198.565 3588.000 200.000 ;
      LAYER met4 ;
        RECT 3483.400 196.955 3588.000 198.165 ;
        RECT 3385.670 176.425 3444.005 176.690 ;
        RECT 3445.135 176.425 3588.000 196.955 ;
        RECT 3385.670 175.165 3588.000 176.425 ;
        RECT 1753.030 174.565 1831.035 175.165 ;
        RECT 2299.965 174.565 2373.035 175.165 ;
        RECT 2841.965 174.565 2915.035 175.165 ;
        RECT 3385.255 174.565 3588.000 175.165 ;
      LAYER met4 ;
        RECT 1284.000 169.515 1753.270 174.165 ;
      LAYER met4 ;
        RECT 1753.670 169.115 1830.330 174.565 ;
      LAYER met4 ;
        RECT 1830.730 169.515 2300.270 174.165 ;
      LAYER met4 ;
        RECT 2300.670 169.115 2372.330 174.565 ;
      LAYER met4 ;
        RECT 2372.730 169.515 2842.270 174.165 ;
      LAYER met4 ;
        RECT 2842.670 169.115 2914.330 174.565 ;
      LAYER met4 ;
        RECT 2914.730 169.515 3385.270 174.165 ;
      LAYER met4 ;
        RECT 3385.670 169.115 3588.000 174.565 ;
        RECT 1753.030 168.515 1831.035 169.115 ;
        RECT 2299.965 168.515 2373.035 169.115 ;
        RECT 2841.965 168.515 2915.035 169.115 ;
        RECT 3385.255 168.515 3588.000 169.115 ;
      LAYER met4 ;
        RECT 1284.000 164.665 1753.270 168.115 ;
      LAYER met4 ;
        RECT 1753.670 164.265 1830.330 168.515 ;
      LAYER met4 ;
        RECT 1830.730 164.665 2300.270 168.115 ;
      LAYER met4 ;
        RECT 2300.670 164.265 2372.330 168.515 ;
      LAYER met4 ;
        RECT 2372.730 164.665 2842.270 168.115 ;
      LAYER met4 ;
        RECT 2842.670 164.265 2914.330 168.515 ;
      LAYER met4 ;
        RECT 2914.730 164.665 3385.270 168.115 ;
      LAYER met4 ;
        RECT 3385.670 164.265 3588.000 168.515 ;
        RECT 1753.030 163.665 1831.035 164.265 ;
        RECT 2299.965 163.665 2373.035 164.265 ;
        RECT 2841.965 163.665 2915.035 164.265 ;
        RECT 3385.255 163.665 3588.000 164.265 ;
      LAYER met4 ;
        RECT 1284.000 159.815 1753.270 163.265 ;
      LAYER met4 ;
        RECT 1753.670 159.415 1830.330 163.665 ;
      LAYER met4 ;
        RECT 1830.730 159.815 2300.270 163.265 ;
      LAYER met4 ;
        RECT 2300.670 159.415 2372.330 163.665 ;
      LAYER met4 ;
        RECT 2372.730 159.815 2842.270 163.265 ;
      LAYER met4 ;
        RECT 2842.670 159.415 2914.330 163.665 ;
      LAYER met4 ;
        RECT 2914.730 159.815 3385.270 163.265 ;
      LAYER met4 ;
        RECT 3385.670 159.415 3588.000 163.665 ;
        RECT 1753.030 158.815 1831.035 159.415 ;
        RECT 2299.965 158.815 2373.035 159.415 ;
        RECT 2841.965 158.815 2915.035 159.415 ;
        RECT 3385.255 158.815 3588.000 159.415 ;
      LAYER met4 ;
        RECT 1284.000 153.765 1753.270 158.415 ;
      LAYER met4 ;
        RECT 1753.670 153.365 1830.330 158.815 ;
      LAYER met4 ;
        RECT 1830.730 153.765 2300.270 158.415 ;
      LAYER met4 ;
        RECT 2300.670 153.365 2372.330 158.815 ;
      LAYER met4 ;
        RECT 2372.730 153.765 2842.270 158.415 ;
      LAYER met4 ;
        RECT 2842.670 153.365 2914.330 158.815 ;
      LAYER met4 ;
        RECT 2914.730 153.765 3385.270 158.415 ;
      LAYER met4 ;
        RECT 3385.670 153.365 3588.000 158.815 ;
        RECT 1753.030 152.665 1831.035 153.365 ;
        RECT 2299.965 152.665 2373.035 153.365 ;
        RECT 2841.965 152.665 2915.035 153.365 ;
        RECT 3385.255 152.665 3588.000 153.365 ;
      LAYER met4 ;
        RECT 1284.000 151.935 1784.910 152.265 ;
      LAYER met4 ;
        RECT 1785.310 152.035 1828.990 152.665 ;
      LAYER met4 ;
        RECT 1829.390 151.935 3407.575 152.265 ;
      LAYER met4 ;
        RECT 0.000 147.275 178.050 148.755 ;
      LAYER met4 ;
        RECT 179.065 148.655 1777.535 151.635 ;
      LAYER met4 ;
        RECT 0.000 143.995 176.690 147.275 ;
      LAYER met4 ;
        RECT 178.450 147.175 200.000 148.355 ;
      LAYER met4 ;
        RECT 200.000 147.275 667.000 148.255 ;
      LAYER met4 ;
        RECT 667.000 147.175 668.270 148.355 ;
      LAYER met4 ;
        RECT 668.670 147.275 740.330 148.255 ;
      LAYER met4 ;
        RECT 740.730 147.175 742.000 148.355 ;
      LAYER met4 ;
        RECT 742.000 147.275 1752.000 148.255 ;
      LAYER met4 ;
        RECT 1752.000 147.175 1753.270 148.355 ;
      LAYER met4 ;
        RECT 1777.935 148.255 1779.455 151.535 ;
      LAYER met4 ;
        RECT 1779.855 148.655 3404.875 151.635 ;
      LAYER met4 ;
        RECT 3407.975 151.535 3588.000 152.665 ;
        RECT 3405.275 148.755 3588.000 151.535 ;
        RECT 1753.670 147.275 1830.330 148.255 ;
        RECT 0.000 142.865 176.425 143.995 ;
      LAYER met4 ;
        RECT 177.090 143.895 1793.240 146.875 ;
        RECT 176.825 143.265 668.270 143.595 ;
      LAYER met4 ;
        RECT 668.670 142.865 740.330 143.495 ;
      LAYER met4 ;
        RECT 740.730 143.265 1209.000 143.595 ;
      LAYER met4 ;
        RECT 1209.000 142.865 1284.000 143.495 ;
      LAYER met4 ;
        RECT 1284.000 143.265 1784.910 143.595 ;
      LAYER met4 ;
        RECT 1793.640 143.495 1795.160 147.275 ;
      LAYER met4 ;
        RECT 1830.730 147.175 1832.000 148.355 ;
      LAYER met4 ;
        RECT 1832.000 147.275 2299.000 148.255 ;
      LAYER met4 ;
        RECT 2299.000 147.175 2300.270 148.355 ;
      LAYER met4 ;
        RECT 2300.670 147.275 2372.330 148.255 ;
      LAYER met4 ;
        RECT 2372.730 147.175 2374.000 148.355 ;
      LAYER met4 ;
        RECT 2374.000 147.275 2841.000 148.255 ;
      LAYER met4 ;
        RECT 2841.000 147.175 2842.270 148.355 ;
      LAYER met4 ;
        RECT 2842.670 147.275 2914.330 148.255 ;
      LAYER met4 ;
        RECT 2914.730 147.175 2916.000 148.355 ;
      LAYER met4 ;
        RECT 2916.000 147.275 3384.000 148.255 ;
      LAYER met4 ;
        RECT 3384.000 147.175 3405.555 148.355 ;
      LAYER met4 ;
        RECT 3405.955 147.275 3588.000 148.755 ;
      LAYER met4 ;
        RECT 1795.560 143.895 3410.910 146.875 ;
      LAYER met4 ;
        RECT 3411.310 143.995 3588.000 147.275 ;
        RECT 1785.310 142.865 1828.990 143.495 ;
      LAYER met4 ;
        RECT 1829.390 143.265 3411.175 143.595 ;
      LAYER met4 ;
        RECT 3411.575 142.865 3588.000 143.995 ;
        RECT 0.000 142.165 667.000 142.865 ;
        RECT 667.965 142.165 741.035 142.865 ;
        RECT 742.000 142.165 1752.000 142.865 ;
        RECT 1753.030 142.165 1831.035 142.865 ;
        RECT 1832.000 142.165 2299.000 142.865 ;
        RECT 2299.965 142.165 2373.035 142.865 ;
        RECT 2374.000 142.165 2841.000 142.865 ;
        RECT 2841.965 142.165 2915.035 142.865 ;
        RECT 2916.000 142.165 3384.000 142.865 ;
        RECT 3385.255 142.165 3588.000 142.865 ;
        RECT 0.000 136.915 197.975 142.165 ;
      LAYER met4 ;
        RECT 198.375 137.315 668.270 141.765 ;
      LAYER met4 ;
        RECT 668.670 136.915 740.330 142.165 ;
      LAYER met4 ;
        RECT 740.730 137.315 1209.000 141.765 ;
      LAYER met4 ;
        RECT 1209.000 136.915 1284.000 142.165 ;
      LAYER met4 ;
        RECT 1284.000 137.315 1753.270 141.765 ;
      LAYER met4 ;
        RECT 1753.670 136.915 1830.330 142.165 ;
      LAYER met4 ;
        RECT 1830.730 137.315 2300.270 141.765 ;
      LAYER met4 ;
        RECT 2300.670 136.915 2372.330 142.165 ;
      LAYER met4 ;
        RECT 2372.730 137.315 2842.270 141.765 ;
      LAYER met4 ;
        RECT 2842.670 136.915 2914.330 142.165 ;
      LAYER met4 ;
        RECT 2914.730 137.315 3385.270 141.765 ;
      LAYER met4 ;
        RECT 3385.670 136.915 3588.000 142.165 ;
        RECT 0.000 136.315 665.000 136.915 ;
        RECT 667.965 136.315 741.035 136.915 ;
        RECT 742.000 136.315 1207.000 136.915 ;
        RECT 1209.000 136.315 1749.000 136.915 ;
        RECT 1753.030 136.315 1831.035 136.915 ;
        RECT 1832.000 136.315 2297.000 136.915 ;
        RECT 2299.965 136.315 2373.035 136.915 ;
        RECT 2374.000 136.315 2839.000 136.915 ;
        RECT 2841.965 136.315 2915.035 136.915 ;
        RECT 2916.000 136.315 3381.000 136.915 ;
        RECT 3385.255 136.315 3588.000 136.915 ;
        RECT 0.000 131.065 198.120 136.315 ;
      LAYER met4 ;
        RECT 198.520 131.465 668.270 135.915 ;
      LAYER met4 ;
        RECT 668.670 131.065 740.330 136.315 ;
      LAYER met4 ;
        RECT 740.730 131.465 1209.000 135.915 ;
      LAYER met4 ;
        RECT 1209.000 131.065 1284.000 136.315 ;
      LAYER met4 ;
        RECT 1284.000 131.465 1753.270 135.915 ;
      LAYER met4 ;
        RECT 1753.670 131.065 1830.330 136.315 ;
      LAYER met4 ;
        RECT 1830.730 131.465 2300.270 135.915 ;
      LAYER met4 ;
        RECT 2300.670 131.065 2372.330 136.315 ;
      LAYER met4 ;
        RECT 2372.730 131.465 2842.270 135.915 ;
      LAYER met4 ;
        RECT 2842.670 131.065 2914.330 136.315 ;
      LAYER met4 ;
        RECT 2914.730 131.465 3385.270 135.915 ;
      LAYER met4 ;
        RECT 3385.670 131.065 3588.000 136.315 ;
        RECT 0.000 130.365 667.000 131.065 ;
        RECT 667.965 130.365 741.035 131.065 ;
        RECT 0.000 104.600 196.955 130.365 ;
        RECT 200.000 129.965 667.000 130.365 ;
      LAYER met4 ;
        RECT 197.355 105.000 201.000 129.965 ;
      LAYER met4 ;
        RECT 201.000 105.000 219.000 129.965 ;
      LAYER met4 ;
        RECT 219.000 105.000 221.000 129.965 ;
      LAYER met4 ;
        RECT 221.000 105.000 239.000 129.965 ;
      LAYER met4 ;
        RECT 239.000 105.000 241.000 129.965 ;
      LAYER met4 ;
        RECT 241.000 105.000 259.000 129.965 ;
      LAYER met4 ;
        RECT 259.000 105.000 261.000 129.965 ;
      LAYER met4 ;
        RECT 261.000 105.000 279.000 129.965 ;
      LAYER met4 ;
        RECT 279.000 105.000 281.000 129.965 ;
      LAYER met4 ;
        RECT 281.000 105.000 299.000 129.965 ;
      LAYER met4 ;
        RECT 299.000 105.000 301.000 129.965 ;
      LAYER met4 ;
        RECT 301.000 105.000 319.000 129.965 ;
      LAYER met4 ;
        RECT 319.000 105.000 321.000 129.965 ;
      LAYER met4 ;
        RECT 321.000 105.000 339.000 129.965 ;
      LAYER met4 ;
        RECT 339.000 105.000 341.000 129.965 ;
      LAYER met4 ;
        RECT 341.000 105.000 359.000 129.965 ;
      LAYER met4 ;
        RECT 359.000 105.000 361.000 129.965 ;
      LAYER met4 ;
        RECT 361.000 105.000 379.000 129.965 ;
      LAYER met4 ;
        RECT 379.000 105.000 381.000 129.965 ;
      LAYER met4 ;
        RECT 381.000 105.000 399.000 129.965 ;
      LAYER met4 ;
        RECT 399.000 105.000 401.000 129.965 ;
      LAYER met4 ;
        RECT 401.000 105.000 419.000 129.965 ;
      LAYER met4 ;
        RECT 419.000 105.000 421.000 129.965 ;
      LAYER met4 ;
        RECT 421.000 105.000 439.000 129.965 ;
      LAYER met4 ;
        RECT 439.000 105.000 441.000 129.965 ;
      LAYER met4 ;
        RECT 441.000 105.000 459.000 129.965 ;
      LAYER met4 ;
        RECT 459.000 105.000 461.000 129.965 ;
      LAYER met4 ;
        RECT 461.000 105.000 479.000 129.965 ;
      LAYER met4 ;
        RECT 479.000 105.000 481.000 129.965 ;
      LAYER met4 ;
        RECT 481.000 105.000 499.000 129.965 ;
      LAYER met4 ;
        RECT 499.000 105.000 501.000 129.965 ;
      LAYER met4 ;
        RECT 501.000 105.000 519.000 129.965 ;
      LAYER met4 ;
        RECT 519.000 105.000 521.000 129.965 ;
      LAYER met4 ;
        RECT 521.000 105.000 539.000 129.965 ;
      LAYER met4 ;
        RECT 539.000 105.000 541.000 129.965 ;
      LAYER met4 ;
        RECT 541.000 105.000 559.000 129.965 ;
      LAYER met4 ;
        RECT 559.000 105.000 561.000 129.965 ;
      LAYER met4 ;
        RECT 561.000 105.000 579.000 129.965 ;
      LAYER met4 ;
        RECT 579.000 105.000 581.000 129.965 ;
      LAYER met4 ;
        RECT 581.000 105.000 599.000 129.965 ;
      LAYER met4 ;
        RECT 599.000 105.000 601.000 129.965 ;
      LAYER met4 ;
        RECT 601.000 105.000 619.000 129.965 ;
      LAYER met4 ;
        RECT 619.000 105.000 621.000 129.965 ;
      LAYER met4 ;
        RECT 621.000 105.000 639.000 129.965 ;
      LAYER met4 ;
        RECT 639.000 105.000 641.000 129.965 ;
      LAYER met4 ;
        RECT 641.000 105.000 659.000 129.965 ;
      LAYER met4 ;
        RECT 659.000 105.000 661.000 129.965 ;
      LAYER met4 ;
        RECT 661.000 105.000 664.000 129.965 ;
      LAYER met4 ;
        RECT 664.000 105.000 668.270 129.965 ;
      LAYER met4 ;
        RECT 200.000 104.600 667.000 105.000 ;
        RECT 668.670 104.600 740.330 130.365 ;
        RECT 742.000 129.965 1752.000 131.065 ;
        RECT 1753.030 130.365 1831.035 131.065 ;
      LAYER met4 ;
        RECT 740.730 105.000 743.000 129.965 ;
      LAYER met4 ;
        RECT 743.000 105.000 761.000 129.965 ;
      LAYER met4 ;
        RECT 761.000 105.000 763.000 129.965 ;
      LAYER met4 ;
        RECT 763.000 105.000 781.000 129.965 ;
      LAYER met4 ;
        RECT 781.000 105.000 783.000 129.965 ;
      LAYER met4 ;
        RECT 783.000 105.000 801.000 129.965 ;
      LAYER met4 ;
        RECT 801.000 105.000 803.000 129.965 ;
      LAYER met4 ;
        RECT 803.000 105.000 821.000 129.965 ;
      LAYER met4 ;
        RECT 821.000 105.000 823.000 129.965 ;
      LAYER met4 ;
        RECT 823.000 105.000 841.000 129.965 ;
      LAYER met4 ;
        RECT 841.000 105.000 843.000 129.965 ;
      LAYER met4 ;
        RECT 843.000 105.000 861.000 129.965 ;
      LAYER met4 ;
        RECT 861.000 105.000 863.000 129.965 ;
      LAYER met4 ;
        RECT 863.000 105.000 881.000 129.965 ;
      LAYER met4 ;
        RECT 881.000 105.000 883.000 129.965 ;
      LAYER met4 ;
        RECT 883.000 105.000 901.000 129.965 ;
      LAYER met4 ;
        RECT 901.000 105.000 903.000 129.965 ;
      LAYER met4 ;
        RECT 903.000 105.000 921.000 129.965 ;
      LAYER met4 ;
        RECT 921.000 105.000 923.000 129.965 ;
      LAYER met4 ;
        RECT 923.000 105.000 941.000 129.965 ;
      LAYER met4 ;
        RECT 941.000 105.000 943.000 129.965 ;
      LAYER met4 ;
        RECT 943.000 105.000 961.000 129.965 ;
      LAYER met4 ;
        RECT 961.000 105.000 963.000 129.965 ;
      LAYER met4 ;
        RECT 963.000 105.000 981.000 129.965 ;
      LAYER met4 ;
        RECT 981.000 105.000 983.000 129.965 ;
      LAYER met4 ;
        RECT 983.000 105.000 1001.000 129.965 ;
      LAYER met4 ;
        RECT 1001.000 105.000 1003.000 129.965 ;
      LAYER met4 ;
        RECT 1003.000 105.000 1021.000 129.965 ;
      LAYER met4 ;
        RECT 1021.000 105.000 1023.000 129.965 ;
      LAYER met4 ;
        RECT 1023.000 105.000 1041.000 129.965 ;
      LAYER met4 ;
        RECT 1041.000 105.000 1043.000 129.965 ;
      LAYER met4 ;
        RECT 1043.000 105.000 1061.000 129.965 ;
      LAYER met4 ;
        RECT 1061.000 105.000 1063.000 129.965 ;
      LAYER met4 ;
        RECT 1063.000 105.000 1081.000 129.965 ;
      LAYER met4 ;
        RECT 1081.000 105.000 1083.000 129.965 ;
      LAYER met4 ;
        RECT 1083.000 105.000 1101.000 129.965 ;
      LAYER met4 ;
        RECT 1101.000 105.000 1103.000 129.965 ;
      LAYER met4 ;
        RECT 1103.000 105.000 1121.000 129.965 ;
      LAYER met4 ;
        RECT 1121.000 105.000 1123.000 129.965 ;
      LAYER met4 ;
        RECT 1123.000 105.000 1141.000 129.965 ;
      LAYER met4 ;
        RECT 1141.000 105.000 1143.000 129.965 ;
      LAYER met4 ;
        RECT 1143.000 105.000 1161.000 129.965 ;
      LAYER met4 ;
        RECT 1161.000 105.000 1163.000 129.965 ;
      LAYER met4 ;
        RECT 1163.000 105.000 1181.000 129.965 ;
      LAYER met4 ;
        RECT 1181.000 105.000 1183.000 129.965 ;
      LAYER met4 ;
        RECT 1183.000 105.000 1201.000 129.965 ;
      LAYER met4 ;
        RECT 1201.000 105.000 1203.000 129.965 ;
      LAYER met4 ;
        RECT 1203.000 105.000 1206.000 129.965 ;
      LAYER met4 ;
        RECT 1206.000 105.000 1209.000 129.965 ;
      LAYER met4 ;
        RECT 1209.000 105.000 1284.000 129.965 ;
      LAYER met4 ;
        RECT 1284.000 105.000 1285.000 129.965 ;
      LAYER met4 ;
        RECT 1285.000 105.000 1303.000 129.965 ;
      LAYER met4 ;
        RECT 1303.000 105.000 1305.000 129.965 ;
      LAYER met4 ;
        RECT 1305.000 105.000 1323.000 129.965 ;
      LAYER met4 ;
        RECT 1323.000 105.000 1325.000 129.965 ;
      LAYER met4 ;
        RECT 1325.000 105.000 1343.000 129.965 ;
      LAYER met4 ;
        RECT 1343.000 105.000 1345.000 129.965 ;
      LAYER met4 ;
        RECT 1345.000 105.000 1363.000 129.965 ;
      LAYER met4 ;
        RECT 1363.000 105.000 1365.000 129.965 ;
      LAYER met4 ;
        RECT 1365.000 105.000 1383.000 129.965 ;
      LAYER met4 ;
        RECT 1383.000 105.000 1385.000 129.965 ;
      LAYER met4 ;
        RECT 1385.000 105.000 1403.000 129.965 ;
      LAYER met4 ;
        RECT 1403.000 105.000 1405.000 129.965 ;
      LAYER met4 ;
        RECT 1405.000 105.000 1423.000 129.965 ;
      LAYER met4 ;
        RECT 1423.000 105.000 1425.000 129.965 ;
      LAYER met4 ;
        RECT 1425.000 105.000 1443.000 129.965 ;
      LAYER met4 ;
        RECT 1443.000 105.000 1445.000 129.965 ;
      LAYER met4 ;
        RECT 1445.000 105.000 1463.000 129.965 ;
      LAYER met4 ;
        RECT 1463.000 105.000 1465.000 129.965 ;
      LAYER met4 ;
        RECT 1465.000 105.000 1483.000 129.965 ;
      LAYER met4 ;
        RECT 1483.000 105.000 1485.000 129.965 ;
      LAYER met4 ;
        RECT 1485.000 105.000 1503.000 129.965 ;
      LAYER met4 ;
        RECT 1503.000 105.000 1505.000 129.965 ;
      LAYER met4 ;
        RECT 1505.000 105.000 1523.000 129.965 ;
      LAYER met4 ;
        RECT 1523.000 105.000 1525.000 129.965 ;
      LAYER met4 ;
        RECT 1525.000 105.000 1543.000 129.965 ;
      LAYER met4 ;
        RECT 1543.000 105.000 1545.000 129.965 ;
      LAYER met4 ;
        RECT 1545.000 105.000 1563.000 129.965 ;
      LAYER met4 ;
        RECT 1563.000 105.000 1565.000 129.965 ;
      LAYER met4 ;
        RECT 1565.000 105.000 1583.000 129.965 ;
      LAYER met4 ;
        RECT 1583.000 105.000 1585.000 129.965 ;
      LAYER met4 ;
        RECT 1585.000 105.000 1603.000 129.965 ;
      LAYER met4 ;
        RECT 1603.000 105.000 1605.000 129.965 ;
      LAYER met4 ;
        RECT 1605.000 105.000 1623.000 129.965 ;
      LAYER met4 ;
        RECT 1623.000 105.000 1625.000 129.965 ;
      LAYER met4 ;
        RECT 1625.000 105.000 1643.000 129.965 ;
      LAYER met4 ;
        RECT 1643.000 105.000 1645.000 129.965 ;
      LAYER met4 ;
        RECT 1645.000 105.000 1663.000 129.965 ;
      LAYER met4 ;
        RECT 1663.000 105.000 1665.000 129.965 ;
      LAYER met4 ;
        RECT 1665.000 105.000 1683.000 129.965 ;
      LAYER met4 ;
        RECT 1683.000 105.000 1685.000 129.965 ;
      LAYER met4 ;
        RECT 1685.000 105.000 1703.000 129.965 ;
      LAYER met4 ;
        RECT 1703.000 105.000 1705.000 129.965 ;
      LAYER met4 ;
        RECT 1705.000 105.000 1723.000 129.965 ;
      LAYER met4 ;
        RECT 1723.000 105.000 1725.000 129.965 ;
      LAYER met4 ;
        RECT 1725.000 105.000 1743.000 129.965 ;
      LAYER met4 ;
        RECT 1743.000 105.000 1745.000 129.965 ;
      LAYER met4 ;
        RECT 1745.000 105.000 1748.000 129.965 ;
      LAYER met4 ;
        RECT 1748.000 105.000 1753.270 129.965 ;
      LAYER met4 ;
        RECT 0.000 102.965 667.000 104.600 ;
        RECT 0.000 25.965 200.000 102.965 ;
        RECT 0.000 24.615 667.000 25.965 ;
        RECT 667.965 24.615 741.035 104.600 ;
        RECT 742.000 102.965 1752.000 105.000 ;
        RECT 1753.670 104.600 1830.330 130.365 ;
        RECT 1832.000 129.965 2299.000 131.065 ;
        RECT 2299.965 130.365 2373.035 131.065 ;
      LAYER met4 ;
        RECT 1830.730 105.000 1833.000 129.965 ;
      LAYER met4 ;
        RECT 1833.000 105.000 1851.000 129.965 ;
      LAYER met4 ;
        RECT 1851.000 105.000 1853.000 129.965 ;
      LAYER met4 ;
        RECT 1853.000 105.000 1871.000 129.965 ;
      LAYER met4 ;
        RECT 1871.000 105.000 1873.000 129.965 ;
      LAYER met4 ;
        RECT 1873.000 105.000 1891.000 129.965 ;
      LAYER met4 ;
        RECT 1891.000 105.000 1893.000 129.965 ;
      LAYER met4 ;
        RECT 1893.000 105.000 1911.000 129.965 ;
      LAYER met4 ;
        RECT 1911.000 105.000 1913.000 129.965 ;
      LAYER met4 ;
        RECT 1913.000 105.000 1931.000 129.965 ;
      LAYER met4 ;
        RECT 1931.000 105.000 1933.000 129.965 ;
      LAYER met4 ;
        RECT 1933.000 105.000 1951.000 129.965 ;
      LAYER met4 ;
        RECT 1951.000 105.000 1953.000 129.965 ;
      LAYER met4 ;
        RECT 1953.000 105.000 1971.000 129.965 ;
      LAYER met4 ;
        RECT 1971.000 105.000 1973.000 129.965 ;
      LAYER met4 ;
        RECT 1973.000 105.000 1991.000 129.965 ;
      LAYER met4 ;
        RECT 1991.000 105.000 1993.000 129.965 ;
      LAYER met4 ;
        RECT 1993.000 105.000 2011.000 129.965 ;
      LAYER met4 ;
        RECT 2011.000 105.000 2013.000 129.965 ;
      LAYER met4 ;
        RECT 2013.000 105.000 2031.000 129.965 ;
      LAYER met4 ;
        RECT 2031.000 105.000 2033.000 129.965 ;
      LAYER met4 ;
        RECT 2033.000 105.000 2051.000 129.965 ;
      LAYER met4 ;
        RECT 2051.000 105.000 2053.000 129.965 ;
      LAYER met4 ;
        RECT 2053.000 105.000 2071.000 129.965 ;
      LAYER met4 ;
        RECT 2071.000 105.000 2073.000 129.965 ;
      LAYER met4 ;
        RECT 2073.000 105.000 2091.000 129.965 ;
      LAYER met4 ;
        RECT 2091.000 105.000 2093.000 129.965 ;
      LAYER met4 ;
        RECT 2093.000 105.000 2111.000 129.965 ;
      LAYER met4 ;
        RECT 2111.000 105.000 2113.000 129.965 ;
      LAYER met4 ;
        RECT 2113.000 105.000 2131.000 129.965 ;
      LAYER met4 ;
        RECT 2131.000 105.000 2133.000 129.965 ;
      LAYER met4 ;
        RECT 2133.000 105.000 2151.000 129.965 ;
      LAYER met4 ;
        RECT 2151.000 105.000 2153.000 129.965 ;
      LAYER met4 ;
        RECT 2153.000 105.000 2171.000 129.965 ;
      LAYER met4 ;
        RECT 2171.000 105.000 2173.000 129.965 ;
      LAYER met4 ;
        RECT 2173.000 105.000 2191.000 129.965 ;
      LAYER met4 ;
        RECT 2191.000 105.000 2193.000 129.965 ;
      LAYER met4 ;
        RECT 2193.000 105.000 2211.000 129.965 ;
      LAYER met4 ;
        RECT 2211.000 105.000 2213.000 129.965 ;
      LAYER met4 ;
        RECT 2213.000 105.000 2231.000 129.965 ;
      LAYER met4 ;
        RECT 2231.000 105.000 2233.000 129.965 ;
      LAYER met4 ;
        RECT 2233.000 105.000 2251.000 129.965 ;
      LAYER met4 ;
        RECT 2251.000 105.000 2253.000 129.965 ;
      LAYER met4 ;
        RECT 2253.000 105.000 2271.000 129.965 ;
      LAYER met4 ;
        RECT 2271.000 105.000 2273.000 129.965 ;
      LAYER met4 ;
        RECT 2273.000 105.000 2291.000 129.965 ;
      LAYER met4 ;
        RECT 2291.000 105.000 2293.000 129.965 ;
      LAYER met4 ;
        RECT 2293.000 105.000 2296.000 129.965 ;
      LAYER met4 ;
        RECT 2296.000 105.000 2300.270 129.965 ;
      LAYER met4 ;
        RECT 1209.000 25.965 1284.000 102.965 ;
        RECT 0.000 0.000 198.165 24.615 ;
      LAYER met4 ;
        RECT 198.565 0.000 200.000 24.215 ;
      LAYER met4 ;
        RECT 200.000 0.000 667.000 24.615 ;
      LAYER met4 ;
        RECT 667.000 0.000 668.270 24.215 ;
      LAYER met4 ;
        RECT 668.670 0.000 740.330 24.615 ;
      LAYER met4 ;
        RECT 740.730 0.000 742.000 24.215 ;
      LAYER met4 ;
        RECT 742.000 0.000 1752.000 25.965 ;
        RECT 1753.030 24.615 1831.035 104.600 ;
        RECT 1832.000 102.965 2299.000 105.000 ;
        RECT 2300.670 104.600 2372.330 130.365 ;
        RECT 2374.000 129.965 2841.000 131.065 ;
        RECT 2841.965 130.365 2915.035 131.065 ;
      LAYER met4 ;
        RECT 2372.730 105.000 2375.000 129.965 ;
      LAYER met4 ;
        RECT 2375.000 105.000 2393.000 129.965 ;
      LAYER met4 ;
        RECT 2393.000 105.000 2395.000 129.965 ;
      LAYER met4 ;
        RECT 2395.000 105.000 2413.000 129.965 ;
      LAYER met4 ;
        RECT 2413.000 105.000 2415.000 129.965 ;
      LAYER met4 ;
        RECT 2415.000 105.000 2433.000 129.965 ;
      LAYER met4 ;
        RECT 2433.000 105.000 2435.000 129.965 ;
      LAYER met4 ;
        RECT 2435.000 105.000 2453.000 129.965 ;
      LAYER met4 ;
        RECT 2453.000 105.000 2455.000 129.965 ;
      LAYER met4 ;
        RECT 2455.000 105.000 2473.000 129.965 ;
      LAYER met4 ;
        RECT 2473.000 105.000 2475.000 129.965 ;
      LAYER met4 ;
        RECT 2475.000 105.000 2493.000 129.965 ;
      LAYER met4 ;
        RECT 2493.000 105.000 2495.000 129.965 ;
      LAYER met4 ;
        RECT 2495.000 105.000 2513.000 129.965 ;
      LAYER met4 ;
        RECT 2513.000 105.000 2515.000 129.965 ;
      LAYER met4 ;
        RECT 2515.000 105.000 2533.000 129.965 ;
      LAYER met4 ;
        RECT 2533.000 105.000 2535.000 129.965 ;
      LAYER met4 ;
        RECT 2535.000 105.000 2553.000 129.965 ;
      LAYER met4 ;
        RECT 2553.000 105.000 2555.000 129.965 ;
      LAYER met4 ;
        RECT 2555.000 105.000 2573.000 129.965 ;
      LAYER met4 ;
        RECT 2573.000 105.000 2575.000 129.965 ;
      LAYER met4 ;
        RECT 2575.000 105.000 2593.000 129.965 ;
      LAYER met4 ;
        RECT 2593.000 105.000 2595.000 129.965 ;
      LAYER met4 ;
        RECT 2595.000 105.000 2613.000 129.965 ;
      LAYER met4 ;
        RECT 2613.000 105.000 2615.000 129.965 ;
      LAYER met4 ;
        RECT 2615.000 105.000 2633.000 129.965 ;
      LAYER met4 ;
        RECT 2633.000 105.000 2635.000 129.965 ;
      LAYER met4 ;
        RECT 2635.000 105.000 2653.000 129.965 ;
      LAYER met4 ;
        RECT 2653.000 105.000 2655.000 129.965 ;
      LAYER met4 ;
        RECT 2655.000 105.000 2673.000 129.965 ;
      LAYER met4 ;
        RECT 2673.000 105.000 2675.000 129.965 ;
      LAYER met4 ;
        RECT 2675.000 105.000 2693.000 129.965 ;
      LAYER met4 ;
        RECT 2693.000 105.000 2695.000 129.965 ;
      LAYER met4 ;
        RECT 2695.000 105.000 2713.000 129.965 ;
      LAYER met4 ;
        RECT 2713.000 105.000 2715.000 129.965 ;
      LAYER met4 ;
        RECT 2715.000 105.000 2733.000 129.965 ;
      LAYER met4 ;
        RECT 2733.000 105.000 2735.000 129.965 ;
      LAYER met4 ;
        RECT 2735.000 105.000 2753.000 129.965 ;
      LAYER met4 ;
        RECT 2753.000 105.000 2755.000 129.965 ;
      LAYER met4 ;
        RECT 2755.000 105.000 2773.000 129.965 ;
      LAYER met4 ;
        RECT 2773.000 105.000 2775.000 129.965 ;
      LAYER met4 ;
        RECT 2775.000 105.000 2793.000 129.965 ;
      LAYER met4 ;
        RECT 2793.000 105.000 2795.000 129.965 ;
      LAYER met4 ;
        RECT 2795.000 105.000 2813.000 129.965 ;
      LAYER met4 ;
        RECT 2813.000 105.000 2815.000 129.965 ;
      LAYER met4 ;
        RECT 2815.000 105.000 2833.000 129.965 ;
      LAYER met4 ;
        RECT 2833.000 105.000 2835.000 129.965 ;
      LAYER met4 ;
        RECT 2835.000 105.000 2838.000 129.965 ;
      LAYER met4 ;
        RECT 2838.000 105.000 2842.270 129.965 ;
        RECT 1752.000 0.000 1753.270 24.215 ;
      LAYER met4 ;
        RECT 1753.670 0.000 1830.330 24.615 ;
      LAYER met4 ;
        RECT 1830.730 0.000 1832.000 24.215 ;
      LAYER met4 ;
        RECT 1832.000 0.000 2299.000 25.965 ;
        RECT 2299.965 24.615 2373.035 104.600 ;
        RECT 2374.000 102.965 2841.000 105.000 ;
        RECT 2842.670 104.600 2914.330 130.365 ;
        RECT 2916.000 129.965 3384.000 131.065 ;
        RECT 3385.255 130.365 3588.000 131.065 ;
      LAYER met4 ;
        RECT 2914.730 105.000 2917.000 129.965 ;
      LAYER met4 ;
        RECT 2917.000 105.000 2935.000 129.965 ;
      LAYER met4 ;
        RECT 2935.000 105.000 2937.000 129.965 ;
      LAYER met4 ;
        RECT 2937.000 105.000 2955.000 129.965 ;
      LAYER met4 ;
        RECT 2955.000 105.000 2957.000 129.965 ;
      LAYER met4 ;
        RECT 2957.000 105.000 2975.000 129.965 ;
      LAYER met4 ;
        RECT 2975.000 105.000 2977.000 129.965 ;
      LAYER met4 ;
        RECT 2977.000 105.000 2995.000 129.965 ;
      LAYER met4 ;
        RECT 2995.000 105.000 2997.000 129.965 ;
      LAYER met4 ;
        RECT 2997.000 105.000 3015.000 129.965 ;
      LAYER met4 ;
        RECT 3015.000 105.000 3017.000 129.965 ;
      LAYER met4 ;
        RECT 3017.000 105.000 3035.000 129.965 ;
      LAYER met4 ;
        RECT 3035.000 105.000 3037.000 129.965 ;
      LAYER met4 ;
        RECT 3037.000 105.000 3055.000 129.965 ;
      LAYER met4 ;
        RECT 3055.000 105.000 3057.000 129.965 ;
      LAYER met4 ;
        RECT 3057.000 105.000 3075.000 129.965 ;
      LAYER met4 ;
        RECT 3075.000 105.000 3077.000 129.965 ;
      LAYER met4 ;
        RECT 3077.000 105.000 3095.000 129.965 ;
      LAYER met4 ;
        RECT 3095.000 105.000 3097.000 129.965 ;
      LAYER met4 ;
        RECT 3097.000 105.000 3115.000 129.965 ;
      LAYER met4 ;
        RECT 3115.000 105.000 3117.000 129.965 ;
      LAYER met4 ;
        RECT 3117.000 105.000 3135.000 129.965 ;
      LAYER met4 ;
        RECT 3135.000 105.000 3137.000 129.965 ;
      LAYER met4 ;
        RECT 3137.000 105.000 3155.000 129.965 ;
      LAYER met4 ;
        RECT 3155.000 105.000 3157.000 129.965 ;
      LAYER met4 ;
        RECT 3157.000 105.000 3175.000 129.965 ;
      LAYER met4 ;
        RECT 3175.000 105.000 3177.000 129.965 ;
      LAYER met4 ;
        RECT 3177.000 105.000 3195.000 129.965 ;
      LAYER met4 ;
        RECT 3195.000 105.000 3197.000 129.965 ;
      LAYER met4 ;
        RECT 3197.000 105.000 3215.000 129.965 ;
      LAYER met4 ;
        RECT 3215.000 105.000 3217.000 129.965 ;
      LAYER met4 ;
        RECT 3217.000 105.000 3235.000 129.965 ;
      LAYER met4 ;
        RECT 3235.000 105.000 3237.000 129.965 ;
      LAYER met4 ;
        RECT 3237.000 105.000 3255.000 129.965 ;
      LAYER met4 ;
        RECT 3255.000 105.000 3257.000 129.965 ;
      LAYER met4 ;
        RECT 3257.000 105.000 3275.000 129.965 ;
      LAYER met4 ;
        RECT 3275.000 105.000 3277.000 129.965 ;
      LAYER met4 ;
        RECT 3277.000 105.000 3295.000 129.965 ;
      LAYER met4 ;
        RECT 3295.000 105.000 3297.000 129.965 ;
      LAYER met4 ;
        RECT 3297.000 105.000 3315.000 129.965 ;
      LAYER met4 ;
        RECT 3315.000 105.000 3317.000 129.965 ;
      LAYER met4 ;
        RECT 3317.000 105.000 3335.000 129.965 ;
      LAYER met4 ;
        RECT 3335.000 105.000 3337.000 129.965 ;
      LAYER met4 ;
        RECT 3337.000 105.000 3355.000 129.965 ;
      LAYER met4 ;
        RECT 3355.000 105.000 3357.000 129.965 ;
      LAYER met4 ;
        RECT 3357.000 105.000 3375.000 129.965 ;
      LAYER met4 ;
        RECT 3375.000 105.000 3377.000 129.965 ;
      LAYER met4 ;
        RECT 3377.000 105.000 3380.000 129.965 ;
      LAYER met4 ;
        RECT 3380.000 105.000 3385.855 129.965 ;
        RECT 2299.000 0.000 2300.270 24.215 ;
      LAYER met4 ;
        RECT 2300.670 0.000 2372.330 24.615 ;
      LAYER met4 ;
        RECT 2372.730 0.000 2374.000 24.215 ;
      LAYER met4 ;
        RECT 2374.000 0.000 2841.000 25.965 ;
        RECT 2841.965 24.615 2915.035 104.600 ;
        RECT 2916.000 102.965 3384.000 105.000 ;
        RECT 3386.255 104.600 3588.000 130.365 ;
      LAYER met4 ;
        RECT 2841.000 0.000 2842.270 24.215 ;
      LAYER met4 ;
        RECT 2842.670 0.000 2914.330 24.615 ;
      LAYER met4 ;
        RECT 2914.730 0.000 2916.000 24.215 ;
      LAYER met4 ;
        RECT 2916.000 0.000 3384.000 25.965 ;
        RECT 3385.255 24.615 3588.000 104.600 ;
      LAYER met4 ;
        RECT 3384.000 0.000 3385.270 24.215 ;
      LAYER met4 ;
        RECT 3385.670 0.000 3588.000 24.615 ;
      LAYER met5 ;
        RECT 0.000 5084.585 204.000 5188.000 ;
      LAYER met5 ;
        RECT 204.000 5163.785 668.000 5188.000 ;
      LAYER met5 ;
        RECT 668.000 5156.610 748.000 5188.000 ;
      LAYER met5 ;
        RECT 748.000 5163.785 1213.000 5188.000 ;
      LAYER met5 ;
        RECT 668.000 5090.960 677.600 5156.610 ;
        RECT 743.400 5090.960 748.000 5156.610 ;
        RECT 668.000 5084.585 748.000 5090.960 ;
        RECT 1213.000 5156.610 1293.000 5188.000 ;
      LAYER met5 ;
        RECT 1293.000 5163.785 1758.000 5188.000 ;
      LAYER met5 ;
        RECT 1213.000 5090.960 1222.600 5156.610 ;
        RECT 1288.400 5090.960 1293.000 5156.610 ;
        RECT 1213.000 5084.585 1293.000 5090.960 ;
        RECT 1758.000 5156.610 1838.000 5188.000 ;
      LAYER met5 ;
        RECT 1838.000 5163.785 2303.000 5188.000 ;
      LAYER met5 ;
        RECT 1758.000 5090.960 1767.600 5156.610 ;
        RECT 1833.400 5090.960 1838.000 5156.610 ;
        RECT 1758.000 5084.585 1838.000 5090.960 ;
        RECT 2303.000 5156.610 2383.000 5188.000 ;
      LAYER met5 ;
        RECT 2383.000 5163.785 2848.000 5188.000 ;
      LAYER met5 ;
        RECT 2303.000 5090.960 2312.600 5156.610 ;
        RECT 2378.400 5090.960 2383.000 5156.610 ;
        RECT 2303.000 5084.585 2383.000 5090.960 ;
        RECT 2848.000 5156.225 2923.000 5188.000 ;
      LAYER met5 ;
        RECT 2923.000 5163.785 3388.000 5188.000 ;
      LAYER met5 ;
        RECT 2848.000 5090.410 2852.500 5156.225 ;
        RECT 2918.400 5090.410 2923.000 5156.225 ;
        RECT 2848.000 5084.585 2923.000 5090.410 ;
        RECT 3388.000 5084.585 3588.000 5188.000 ;
        RECT 0.000 5056.435 200.545 5084.585 ;
      LAYER met5 ;
        RECT 202.145 5058.035 205.000 5082.985 ;
      LAYER met5 ;
        RECT 206.600 5058.035 221.400 5082.985 ;
      LAYER met5 ;
        RECT 223.000 5058.035 225.000 5082.985 ;
      LAYER met5 ;
        RECT 226.600 5058.035 241.400 5082.985 ;
      LAYER met5 ;
        RECT 243.000 5058.035 245.000 5082.985 ;
      LAYER met5 ;
        RECT 246.600 5058.035 261.400 5082.985 ;
      LAYER met5 ;
        RECT 263.000 5058.035 265.000 5082.985 ;
      LAYER met5 ;
        RECT 266.600 5058.035 281.400 5082.985 ;
      LAYER met5 ;
        RECT 283.000 5058.035 285.000 5082.985 ;
      LAYER met5 ;
        RECT 286.600 5058.035 301.400 5082.985 ;
      LAYER met5 ;
        RECT 303.000 5058.035 305.000 5082.985 ;
      LAYER met5 ;
        RECT 306.600 5058.035 321.400 5082.985 ;
      LAYER met5 ;
        RECT 323.000 5058.035 325.000 5082.985 ;
      LAYER met5 ;
        RECT 326.600 5058.035 341.400 5082.985 ;
      LAYER met5 ;
        RECT 343.000 5058.035 345.000 5082.985 ;
      LAYER met5 ;
        RECT 346.600 5058.035 361.400 5082.985 ;
      LAYER met5 ;
        RECT 363.000 5058.035 365.000 5082.985 ;
      LAYER met5 ;
        RECT 366.600 5058.035 381.400 5082.985 ;
      LAYER met5 ;
        RECT 383.000 5058.035 385.000 5082.985 ;
      LAYER met5 ;
        RECT 386.600 5058.035 401.400 5082.985 ;
      LAYER met5 ;
        RECT 403.000 5058.035 405.000 5082.985 ;
      LAYER met5 ;
        RECT 406.600 5058.035 421.400 5082.985 ;
      LAYER met5 ;
        RECT 423.000 5058.035 425.000 5082.985 ;
      LAYER met5 ;
        RECT 426.600 5058.035 441.400 5082.985 ;
      LAYER met5 ;
        RECT 443.000 5058.035 445.000 5082.985 ;
      LAYER met5 ;
        RECT 446.600 5058.035 461.400 5082.985 ;
      LAYER met5 ;
        RECT 463.000 5058.035 465.000 5082.985 ;
      LAYER met5 ;
        RECT 466.600 5058.035 481.400 5082.985 ;
      LAYER met5 ;
        RECT 483.000 5058.035 485.000 5082.985 ;
      LAYER met5 ;
        RECT 486.600 5058.035 501.400 5082.985 ;
      LAYER met5 ;
        RECT 503.000 5058.035 505.000 5082.985 ;
      LAYER met5 ;
        RECT 506.600 5058.035 521.400 5082.985 ;
      LAYER met5 ;
        RECT 523.000 5058.035 525.000 5082.985 ;
      LAYER met5 ;
        RECT 526.600 5058.035 541.400 5082.985 ;
      LAYER met5 ;
        RECT 543.000 5058.035 545.000 5082.985 ;
      LAYER met5 ;
        RECT 546.600 5058.035 561.400 5082.985 ;
      LAYER met5 ;
        RECT 563.000 5058.035 565.000 5082.985 ;
      LAYER met5 ;
        RECT 566.600 5058.035 581.400 5082.985 ;
      LAYER met5 ;
        RECT 583.000 5058.035 585.000 5082.985 ;
      LAYER met5 ;
        RECT 586.600 5058.035 601.400 5082.985 ;
      LAYER met5 ;
        RECT 603.000 5058.035 605.000 5082.985 ;
      LAYER met5 ;
        RECT 606.600 5058.035 621.400 5082.985 ;
      LAYER met5 ;
        RECT 623.000 5058.035 625.000 5082.985 ;
      LAYER met5 ;
        RECT 626.600 5058.035 641.400 5082.985 ;
      LAYER met5 ;
        RECT 643.000 5058.035 645.000 5082.985 ;
      LAYER met5 ;
        RECT 646.600 5058.035 661.400 5082.985 ;
      LAYER met5 ;
        RECT 663.000 5058.035 669.270 5082.985 ;
      LAYER met5 ;
        RECT 0.000 5046.335 201.130 5056.435 ;
      LAYER met5 ;
        RECT 202.730 5052.185 669.270 5056.435 ;
        RECT 202.730 5046.335 669.270 5050.585 ;
      LAYER met5 ;
        RECT 0.000 5034.135 175.245 5046.335 ;
      LAYER met5 ;
        RECT 176.845 5035.735 669.270 5044.735 ;
      LAYER met5 ;
        RECT 0.000 5012.755 201.130 5034.135 ;
      LAYER met5 ;
        RECT 202.730 5029.685 669.270 5034.135 ;
        RECT 202.730 5024.840 669.270 5028.085 ;
        RECT 204.000 5024.835 668.000 5024.840 ;
        RECT 202.730 5019.985 669.270 5023.235 ;
        RECT 202.730 5013.935 669.270 5018.385 ;
      LAYER met5 ;
        RECT 0.000 4992.245 141.665 5012.755 ;
        RECT 0.000 4988.000 103.415 4992.245 ;
        RECT 131.565 4991.225 141.665 4992.245 ;
        RECT 131.565 4991.080 135.815 4991.225 ;
      LAYER met5 ;
        RECT 0.000 4459.000 24.215 4988.000 ;
        RECT 105.015 4983.000 129.965 4990.645 ;
        RECT 105.015 4978.000 129.965 4980.000 ;
      LAYER met5 ;
        RECT 105.015 4961.600 129.965 4976.400 ;
      LAYER met5 ;
        RECT 105.015 4958.000 129.965 4960.000 ;
      LAYER met5 ;
        RECT 105.015 4941.600 129.965 4956.400 ;
      LAYER met5 ;
        RECT 105.015 4938.000 129.965 4940.000 ;
      LAYER met5 ;
        RECT 105.015 4921.600 129.965 4936.400 ;
      LAYER met5 ;
        RECT 105.015 4918.000 129.965 4920.000 ;
      LAYER met5 ;
        RECT 105.015 4901.600 129.965 4916.400 ;
      LAYER met5 ;
        RECT 105.015 4898.000 129.965 4900.000 ;
      LAYER met5 ;
        RECT 105.015 4881.600 129.965 4896.400 ;
      LAYER met5 ;
        RECT 105.015 4878.000 129.965 4880.000 ;
      LAYER met5 ;
        RECT 105.015 4861.600 129.965 4876.400 ;
      LAYER met5 ;
        RECT 105.015 4858.000 129.965 4860.000 ;
      LAYER met5 ;
        RECT 105.015 4841.600 129.965 4856.400 ;
      LAYER met5 ;
        RECT 105.015 4838.000 129.965 4840.000 ;
      LAYER met5 ;
        RECT 105.015 4821.600 129.965 4836.400 ;
      LAYER met5 ;
        RECT 105.015 4818.000 129.965 4820.000 ;
      LAYER met5 ;
        RECT 105.015 4801.600 129.965 4816.400 ;
      LAYER met5 ;
        RECT 105.015 4798.000 129.965 4800.000 ;
      LAYER met5 ;
        RECT 105.015 4781.600 129.965 4796.400 ;
      LAYER met5 ;
        RECT 105.015 4778.000 129.965 4780.000 ;
      LAYER met5 ;
        RECT 105.015 4761.600 129.965 4776.400 ;
      LAYER met5 ;
        RECT 105.015 4758.000 129.965 4760.000 ;
      LAYER met5 ;
        RECT 105.015 4741.600 129.965 4756.400 ;
      LAYER met5 ;
        RECT 105.015 4738.000 129.965 4740.000 ;
      LAYER met5 ;
        RECT 105.015 4721.600 129.965 4736.400 ;
      LAYER met5 ;
        RECT 105.015 4718.000 129.965 4720.000 ;
      LAYER met5 ;
        RECT 105.015 4701.600 129.965 4716.400 ;
      LAYER met5 ;
        RECT 105.015 4698.000 129.965 4700.000 ;
      LAYER met5 ;
        RECT 105.015 4681.600 129.965 4696.400 ;
      LAYER met5 ;
        RECT 105.015 4678.000 129.965 4680.000 ;
      LAYER met5 ;
        RECT 105.015 4661.600 129.965 4676.400 ;
      LAYER met5 ;
        RECT 105.015 4658.000 129.965 4660.000 ;
      LAYER met5 ;
        RECT 105.015 4641.600 129.965 4656.400 ;
      LAYER met5 ;
        RECT 105.015 4638.000 129.965 4640.000 ;
      LAYER met5 ;
        RECT 105.015 4621.600 129.965 4636.400 ;
      LAYER met5 ;
        RECT 105.015 4618.000 129.965 4620.000 ;
      LAYER met5 ;
        RECT 105.015 4601.600 129.965 4616.400 ;
      LAYER met5 ;
        RECT 105.015 4598.000 129.965 4600.000 ;
      LAYER met5 ;
        RECT 105.015 4581.600 129.965 4596.400 ;
      LAYER met5 ;
        RECT 105.015 4578.000 129.965 4580.000 ;
      LAYER met5 ;
        RECT 105.015 4561.600 129.965 4576.400 ;
      LAYER met5 ;
        RECT 105.015 4558.000 129.965 4560.000 ;
      LAYER met5 ;
        RECT 105.015 4541.600 129.965 4556.400 ;
      LAYER met5 ;
        RECT 105.015 4538.000 129.965 4540.000 ;
      LAYER met5 ;
        RECT 105.015 4521.600 129.965 4536.400 ;
      LAYER met5 ;
        RECT 105.015 4518.000 129.965 4520.000 ;
      LAYER met5 ;
        RECT 105.015 4501.600 129.965 4516.400 ;
      LAYER met5 ;
        RECT 105.015 4498.000 129.965 4500.000 ;
      LAYER met5 ;
        RECT 105.015 4481.600 129.965 4496.400 ;
      LAYER met5 ;
        RECT 105.015 4478.000 129.965 4480.000 ;
      LAYER met5 ;
        RECT 105.015 4461.600 129.965 4476.400 ;
        RECT 0.000 4456.130 103.415 4459.000 ;
      LAYER met5 ;
        RECT 105.015 4457.730 129.965 4460.000 ;
        RECT 131.565 4457.730 135.815 4989.480 ;
        RECT 137.415 4457.730 141.665 4989.625 ;
        RECT 143.265 4457.730 152.265 5011.155 ;
      LAYER met5 ;
        RECT 153.865 5006.285 201.130 5012.755 ;
      LAYER met5 ;
        RECT 202.730 5007.885 669.270 5012.335 ;
      LAYER met5 ;
        RECT 670.870 5006.285 745.130 5084.585 ;
      LAYER met5 ;
        RECT 746.730 5058.035 749.000 5082.985 ;
      LAYER met5 ;
        RECT 750.600 5058.035 765.400 5082.985 ;
      LAYER met5 ;
        RECT 767.000 5058.035 769.000 5082.985 ;
      LAYER met5 ;
        RECT 770.600 5058.035 785.400 5082.985 ;
      LAYER met5 ;
        RECT 787.000 5058.035 789.000 5082.985 ;
      LAYER met5 ;
        RECT 790.600 5058.035 805.400 5082.985 ;
      LAYER met5 ;
        RECT 807.000 5058.035 809.000 5082.985 ;
      LAYER met5 ;
        RECT 810.600 5058.035 825.400 5082.985 ;
      LAYER met5 ;
        RECT 827.000 5058.035 829.000 5082.985 ;
      LAYER met5 ;
        RECT 830.600 5058.035 845.400 5082.985 ;
      LAYER met5 ;
        RECT 847.000 5058.035 849.000 5082.985 ;
      LAYER met5 ;
        RECT 850.600 5058.035 865.400 5082.985 ;
      LAYER met5 ;
        RECT 867.000 5058.035 869.000 5082.985 ;
      LAYER met5 ;
        RECT 870.600 5058.035 885.400 5082.985 ;
      LAYER met5 ;
        RECT 887.000 5058.035 889.000 5082.985 ;
      LAYER met5 ;
        RECT 890.600 5058.035 905.400 5082.985 ;
      LAYER met5 ;
        RECT 907.000 5058.035 909.000 5082.985 ;
      LAYER met5 ;
        RECT 910.600 5058.035 925.400 5082.985 ;
      LAYER met5 ;
        RECT 927.000 5058.035 929.000 5082.985 ;
      LAYER met5 ;
        RECT 930.600 5058.035 945.400 5082.985 ;
      LAYER met5 ;
        RECT 947.000 5058.035 949.000 5082.985 ;
      LAYER met5 ;
        RECT 950.600 5058.035 965.400 5082.985 ;
      LAYER met5 ;
        RECT 967.000 5058.035 969.000 5082.985 ;
      LAYER met5 ;
        RECT 970.600 5058.035 985.400 5082.985 ;
      LAYER met5 ;
        RECT 987.000 5058.035 989.000 5082.985 ;
      LAYER met5 ;
        RECT 990.600 5058.035 1005.400 5082.985 ;
      LAYER met5 ;
        RECT 1007.000 5058.035 1009.000 5082.985 ;
      LAYER met5 ;
        RECT 1010.600 5058.035 1025.400 5082.985 ;
      LAYER met5 ;
        RECT 1027.000 5058.035 1029.000 5082.985 ;
      LAYER met5 ;
        RECT 1030.600 5058.035 1045.400 5082.985 ;
      LAYER met5 ;
        RECT 1047.000 5058.035 1049.000 5082.985 ;
      LAYER met5 ;
        RECT 1050.600 5058.035 1065.400 5082.985 ;
      LAYER met5 ;
        RECT 1067.000 5058.035 1069.000 5082.985 ;
      LAYER met5 ;
        RECT 1070.600 5058.035 1085.400 5082.985 ;
      LAYER met5 ;
        RECT 1087.000 5058.035 1089.000 5082.985 ;
      LAYER met5 ;
        RECT 1090.600 5058.035 1105.400 5082.985 ;
      LAYER met5 ;
        RECT 1107.000 5058.035 1109.000 5082.985 ;
      LAYER met5 ;
        RECT 1110.600 5058.035 1125.400 5082.985 ;
      LAYER met5 ;
        RECT 1127.000 5058.035 1129.000 5082.985 ;
      LAYER met5 ;
        RECT 1130.600 5058.035 1145.400 5082.985 ;
      LAYER met5 ;
        RECT 1147.000 5058.035 1149.000 5082.985 ;
      LAYER met5 ;
        RECT 1150.600 5058.035 1165.400 5082.985 ;
      LAYER met5 ;
        RECT 1167.000 5058.035 1169.000 5082.985 ;
      LAYER met5 ;
        RECT 1170.600 5058.035 1185.400 5082.985 ;
      LAYER met5 ;
        RECT 1187.000 5058.035 1189.000 5082.985 ;
      LAYER met5 ;
        RECT 1190.600 5058.035 1205.400 5082.985 ;
      LAYER met5 ;
        RECT 1207.000 5058.035 1209.000 5082.985 ;
        RECT 1212.000 5058.035 1214.270 5082.985 ;
        RECT 746.730 5052.185 1214.270 5056.435 ;
        RECT 746.730 5046.335 1214.270 5050.585 ;
        RECT 746.730 5035.735 1214.270 5044.735 ;
        RECT 746.730 5029.685 1214.270 5034.135 ;
        RECT 746.730 5024.840 1214.270 5028.085 ;
        RECT 748.000 5024.835 1213.000 5024.840 ;
        RECT 746.730 5019.985 1214.270 5023.235 ;
        RECT 746.730 5013.935 1214.270 5018.385 ;
        RECT 746.730 5007.885 1214.270 5012.335 ;
      LAYER met5 ;
        RECT 1215.870 5006.285 1290.130 5084.585 ;
      LAYER met5 ;
        RECT 1291.730 5058.035 1294.000 5082.985 ;
      LAYER met5 ;
        RECT 1295.600 5058.035 1310.400 5082.985 ;
      LAYER met5 ;
        RECT 1312.000 5058.035 1314.000 5082.985 ;
      LAYER met5 ;
        RECT 1315.600 5058.035 1330.400 5082.985 ;
      LAYER met5 ;
        RECT 1332.000 5058.035 1334.000 5082.985 ;
      LAYER met5 ;
        RECT 1335.600 5058.035 1350.400 5082.985 ;
      LAYER met5 ;
        RECT 1352.000 5058.035 1354.000 5082.985 ;
      LAYER met5 ;
        RECT 1355.600 5058.035 1370.400 5082.985 ;
      LAYER met5 ;
        RECT 1372.000 5058.035 1374.000 5082.985 ;
      LAYER met5 ;
        RECT 1375.600 5058.035 1390.400 5082.985 ;
      LAYER met5 ;
        RECT 1392.000 5058.035 1394.000 5082.985 ;
      LAYER met5 ;
        RECT 1395.600 5058.035 1410.400 5082.985 ;
      LAYER met5 ;
        RECT 1412.000 5058.035 1414.000 5082.985 ;
      LAYER met5 ;
        RECT 1415.600 5058.035 1430.400 5082.985 ;
      LAYER met5 ;
        RECT 1432.000 5058.035 1434.000 5082.985 ;
      LAYER met5 ;
        RECT 1435.600 5058.035 1450.400 5082.985 ;
      LAYER met5 ;
        RECT 1452.000 5058.035 1454.000 5082.985 ;
      LAYER met5 ;
        RECT 1455.600 5058.035 1470.400 5082.985 ;
      LAYER met5 ;
        RECT 1472.000 5058.035 1474.000 5082.985 ;
      LAYER met5 ;
        RECT 1475.600 5058.035 1490.400 5082.985 ;
      LAYER met5 ;
        RECT 1492.000 5058.035 1494.000 5082.985 ;
      LAYER met5 ;
        RECT 1495.600 5058.035 1510.400 5082.985 ;
      LAYER met5 ;
        RECT 1512.000 5058.035 1514.000 5082.985 ;
      LAYER met5 ;
        RECT 1515.600 5058.035 1530.400 5082.985 ;
      LAYER met5 ;
        RECT 1532.000 5058.035 1534.000 5082.985 ;
      LAYER met5 ;
        RECT 1535.600 5058.035 1550.400 5082.985 ;
      LAYER met5 ;
        RECT 1552.000 5058.035 1554.000 5082.985 ;
      LAYER met5 ;
        RECT 1555.600 5058.035 1570.400 5082.985 ;
      LAYER met5 ;
        RECT 1572.000 5058.035 1574.000 5082.985 ;
      LAYER met5 ;
        RECT 1575.600 5058.035 1590.400 5082.985 ;
      LAYER met5 ;
        RECT 1592.000 5058.035 1594.000 5082.985 ;
      LAYER met5 ;
        RECT 1595.600 5058.035 1610.400 5082.985 ;
      LAYER met5 ;
        RECT 1612.000 5058.035 1614.000 5082.985 ;
      LAYER met5 ;
        RECT 1615.600 5058.035 1630.400 5082.985 ;
      LAYER met5 ;
        RECT 1632.000 5058.035 1634.000 5082.985 ;
      LAYER met5 ;
        RECT 1635.600 5058.035 1650.400 5082.985 ;
      LAYER met5 ;
        RECT 1652.000 5058.035 1654.000 5082.985 ;
      LAYER met5 ;
        RECT 1655.600 5058.035 1670.400 5082.985 ;
      LAYER met5 ;
        RECT 1672.000 5058.035 1674.000 5082.985 ;
      LAYER met5 ;
        RECT 1675.600 5058.035 1690.400 5082.985 ;
      LAYER met5 ;
        RECT 1692.000 5058.035 1694.000 5082.985 ;
      LAYER met5 ;
        RECT 1695.600 5058.035 1710.400 5082.985 ;
      LAYER met5 ;
        RECT 1712.000 5058.035 1714.000 5082.985 ;
      LAYER met5 ;
        RECT 1715.600 5058.035 1730.400 5082.985 ;
      LAYER met5 ;
        RECT 1732.000 5058.035 1734.000 5082.985 ;
      LAYER met5 ;
        RECT 1735.600 5058.035 1750.400 5082.985 ;
      LAYER met5 ;
        RECT 1752.000 5058.035 1754.000 5082.985 ;
        RECT 1757.000 5058.035 1759.270 5082.985 ;
        RECT 1291.730 5052.185 1759.270 5056.435 ;
        RECT 1291.730 5046.335 1759.270 5050.585 ;
        RECT 1291.730 5035.735 1759.270 5044.735 ;
        RECT 1291.730 5029.685 1759.270 5034.135 ;
        RECT 1291.730 5024.840 1759.270 5028.085 ;
        RECT 1293.000 5024.835 1758.000 5024.840 ;
        RECT 1291.730 5019.985 1759.270 5023.235 ;
        RECT 1291.730 5013.935 1759.270 5018.385 ;
        RECT 1291.730 5007.885 1759.270 5012.335 ;
      LAYER met5 ;
        RECT 1760.870 5006.285 1835.130 5084.585 ;
      LAYER met5 ;
        RECT 1836.730 5058.035 1839.000 5082.985 ;
      LAYER met5 ;
        RECT 1840.600 5058.035 1855.400 5082.985 ;
      LAYER met5 ;
        RECT 1857.000 5058.035 1859.000 5082.985 ;
      LAYER met5 ;
        RECT 1860.600 5058.035 1875.400 5082.985 ;
      LAYER met5 ;
        RECT 1877.000 5058.035 1879.000 5082.985 ;
      LAYER met5 ;
        RECT 1880.600 5058.035 1895.400 5082.985 ;
      LAYER met5 ;
        RECT 1897.000 5058.035 1899.000 5082.985 ;
      LAYER met5 ;
        RECT 1900.600 5058.035 1915.400 5082.985 ;
      LAYER met5 ;
        RECT 1917.000 5058.035 1919.000 5082.985 ;
      LAYER met5 ;
        RECT 1920.600 5058.035 1935.400 5082.985 ;
      LAYER met5 ;
        RECT 1937.000 5058.035 1939.000 5082.985 ;
      LAYER met5 ;
        RECT 1940.600 5058.035 1955.400 5082.985 ;
      LAYER met5 ;
        RECT 1957.000 5058.035 1959.000 5082.985 ;
      LAYER met5 ;
        RECT 1960.600 5058.035 1975.400 5082.985 ;
      LAYER met5 ;
        RECT 1977.000 5058.035 1979.000 5082.985 ;
      LAYER met5 ;
        RECT 1980.600 5058.035 1995.400 5082.985 ;
      LAYER met5 ;
        RECT 1997.000 5058.035 1999.000 5082.985 ;
      LAYER met5 ;
        RECT 2000.600 5058.035 2015.400 5082.985 ;
      LAYER met5 ;
        RECT 2017.000 5058.035 2019.000 5082.985 ;
      LAYER met5 ;
        RECT 2020.600 5058.035 2035.400 5082.985 ;
      LAYER met5 ;
        RECT 2037.000 5058.035 2039.000 5082.985 ;
      LAYER met5 ;
        RECT 2040.600 5058.035 2055.400 5082.985 ;
      LAYER met5 ;
        RECT 2057.000 5058.035 2059.000 5082.985 ;
      LAYER met5 ;
        RECT 2060.600 5058.035 2075.400 5082.985 ;
      LAYER met5 ;
        RECT 2077.000 5058.035 2079.000 5082.985 ;
      LAYER met5 ;
        RECT 2080.600 5058.035 2095.400 5082.985 ;
      LAYER met5 ;
        RECT 2097.000 5058.035 2099.000 5082.985 ;
      LAYER met5 ;
        RECT 2100.600 5058.035 2115.400 5082.985 ;
      LAYER met5 ;
        RECT 2117.000 5058.035 2119.000 5082.985 ;
      LAYER met5 ;
        RECT 2120.600 5058.035 2135.400 5082.985 ;
      LAYER met5 ;
        RECT 2137.000 5058.035 2139.000 5082.985 ;
      LAYER met5 ;
        RECT 2140.600 5058.035 2155.400 5082.985 ;
      LAYER met5 ;
        RECT 2157.000 5058.035 2159.000 5082.985 ;
      LAYER met5 ;
        RECT 2160.600 5058.035 2175.400 5082.985 ;
      LAYER met5 ;
        RECT 2177.000 5058.035 2179.000 5082.985 ;
      LAYER met5 ;
        RECT 2180.600 5058.035 2195.400 5082.985 ;
      LAYER met5 ;
        RECT 2197.000 5058.035 2199.000 5082.985 ;
      LAYER met5 ;
        RECT 2200.600 5058.035 2215.400 5082.985 ;
      LAYER met5 ;
        RECT 2217.000 5058.035 2219.000 5082.985 ;
      LAYER met5 ;
        RECT 2220.600 5058.035 2235.400 5082.985 ;
      LAYER met5 ;
        RECT 2237.000 5058.035 2239.000 5082.985 ;
      LAYER met5 ;
        RECT 2240.600 5058.035 2255.400 5082.985 ;
      LAYER met5 ;
        RECT 2257.000 5058.035 2259.000 5082.985 ;
      LAYER met5 ;
        RECT 2260.600 5058.035 2275.400 5082.985 ;
      LAYER met5 ;
        RECT 2277.000 5058.035 2279.000 5082.985 ;
      LAYER met5 ;
        RECT 2280.600 5058.035 2295.400 5082.985 ;
      LAYER met5 ;
        RECT 2297.000 5058.035 2299.000 5082.985 ;
        RECT 2302.000 5058.035 2304.270 5082.985 ;
        RECT 1836.730 5052.185 2304.270 5056.435 ;
        RECT 1836.730 5046.335 2304.270 5050.585 ;
        RECT 1836.730 5035.735 2304.270 5044.735 ;
        RECT 1836.730 5029.685 2304.270 5034.135 ;
        RECT 1836.730 5024.840 2304.270 5028.085 ;
        RECT 1838.000 5024.835 2303.000 5024.840 ;
        RECT 1836.730 5019.985 2304.270 5023.235 ;
        RECT 1836.730 5013.935 2304.270 5018.385 ;
        RECT 1836.730 5007.885 2304.270 5012.335 ;
      LAYER met5 ;
        RECT 2305.870 5006.285 2380.130 5084.585 ;
      LAYER met5 ;
        RECT 2381.730 5058.035 2384.000 5082.985 ;
      LAYER met5 ;
        RECT 2385.600 5058.035 2400.400 5082.985 ;
      LAYER met5 ;
        RECT 2402.000 5058.035 2404.000 5082.985 ;
      LAYER met5 ;
        RECT 2405.600 5058.035 2420.400 5082.985 ;
      LAYER met5 ;
        RECT 2422.000 5058.035 2424.000 5082.985 ;
      LAYER met5 ;
        RECT 2425.600 5058.035 2440.400 5082.985 ;
      LAYER met5 ;
        RECT 2442.000 5058.035 2444.000 5082.985 ;
      LAYER met5 ;
        RECT 2445.600 5058.035 2460.400 5082.985 ;
      LAYER met5 ;
        RECT 2462.000 5058.035 2464.000 5082.985 ;
      LAYER met5 ;
        RECT 2465.600 5058.035 2480.400 5082.985 ;
      LAYER met5 ;
        RECT 2482.000 5058.035 2484.000 5082.985 ;
      LAYER met5 ;
        RECT 2485.600 5058.035 2500.400 5082.985 ;
      LAYER met5 ;
        RECT 2502.000 5058.035 2504.000 5082.985 ;
      LAYER met5 ;
        RECT 2505.600 5058.035 2520.400 5082.985 ;
      LAYER met5 ;
        RECT 2522.000 5058.035 2524.000 5082.985 ;
      LAYER met5 ;
        RECT 2525.600 5058.035 2540.400 5082.985 ;
      LAYER met5 ;
        RECT 2542.000 5058.035 2544.000 5082.985 ;
      LAYER met5 ;
        RECT 2545.600 5058.035 2560.400 5082.985 ;
      LAYER met5 ;
        RECT 2562.000 5058.035 2564.000 5082.985 ;
      LAYER met5 ;
        RECT 2565.600 5058.035 2580.400 5082.985 ;
      LAYER met5 ;
        RECT 2582.000 5058.035 2584.000 5082.985 ;
      LAYER met5 ;
        RECT 2585.600 5058.035 2600.400 5082.985 ;
      LAYER met5 ;
        RECT 2602.000 5058.035 2604.000 5082.985 ;
      LAYER met5 ;
        RECT 2605.600 5058.035 2620.400 5082.985 ;
      LAYER met5 ;
        RECT 2622.000 5058.035 2624.000 5082.985 ;
      LAYER met5 ;
        RECT 2625.600 5058.035 2640.400 5082.985 ;
      LAYER met5 ;
        RECT 2642.000 5058.035 2644.000 5082.985 ;
      LAYER met5 ;
        RECT 2645.600 5058.035 2660.400 5082.985 ;
      LAYER met5 ;
        RECT 2662.000 5058.035 2664.000 5082.985 ;
      LAYER met5 ;
        RECT 2665.600 5058.035 2680.400 5082.985 ;
      LAYER met5 ;
        RECT 2682.000 5058.035 2684.000 5082.985 ;
      LAYER met5 ;
        RECT 2685.600 5058.035 2700.400 5082.985 ;
      LAYER met5 ;
        RECT 2702.000 5058.035 2704.000 5082.985 ;
      LAYER met5 ;
        RECT 2705.600 5058.035 2720.400 5082.985 ;
      LAYER met5 ;
        RECT 2722.000 5058.035 2724.000 5082.985 ;
      LAYER met5 ;
        RECT 2725.600 5058.035 2740.400 5082.985 ;
      LAYER met5 ;
        RECT 2742.000 5058.035 2744.000 5082.985 ;
      LAYER met5 ;
        RECT 2745.600 5058.035 2760.400 5082.985 ;
      LAYER met5 ;
        RECT 2762.000 5058.035 2764.000 5082.985 ;
      LAYER met5 ;
        RECT 2765.600 5058.035 2780.400 5082.985 ;
      LAYER met5 ;
        RECT 2782.000 5058.035 2784.000 5082.985 ;
      LAYER met5 ;
        RECT 2785.600 5058.035 2800.400 5082.985 ;
      LAYER met5 ;
        RECT 2802.000 5058.035 2804.000 5082.985 ;
      LAYER met5 ;
        RECT 2805.600 5058.035 2820.400 5082.985 ;
      LAYER met5 ;
        RECT 2822.000 5058.035 2824.000 5082.985 ;
      LAYER met5 ;
        RECT 2825.600 5058.035 2840.400 5082.985 ;
      LAYER met5 ;
        RECT 2842.000 5058.035 2844.000 5082.985 ;
        RECT 2847.000 5058.035 2849.270 5082.985 ;
        RECT 2381.730 5052.185 2849.270 5056.435 ;
        RECT 2381.730 5046.335 2849.270 5050.585 ;
        RECT 2381.730 5035.735 2849.270 5044.735 ;
        RECT 2381.730 5029.685 2849.270 5034.135 ;
        RECT 2381.730 5024.840 2849.270 5028.085 ;
        RECT 2383.000 5024.835 2848.000 5024.840 ;
        RECT 2381.730 5019.985 2849.270 5023.235 ;
        RECT 2381.730 5013.935 2849.270 5018.385 ;
        RECT 2381.730 5007.885 2849.270 5012.335 ;
      LAYER met5 ;
        RECT 2850.870 5006.285 2920.130 5084.585 ;
      LAYER met5 ;
        RECT 2921.730 5058.035 2924.000 5082.985 ;
      LAYER met5 ;
        RECT 2925.600 5058.035 2940.400 5082.985 ;
      LAYER met5 ;
        RECT 2942.000 5058.035 2944.000 5082.985 ;
      LAYER met5 ;
        RECT 2945.600 5058.035 2960.400 5082.985 ;
      LAYER met5 ;
        RECT 2962.000 5058.035 2964.000 5082.985 ;
      LAYER met5 ;
        RECT 2965.600 5058.035 2980.400 5082.985 ;
      LAYER met5 ;
        RECT 2982.000 5058.035 2984.000 5082.985 ;
      LAYER met5 ;
        RECT 2985.600 5058.035 3000.400 5082.985 ;
      LAYER met5 ;
        RECT 3002.000 5058.035 3004.000 5082.985 ;
      LAYER met5 ;
        RECT 3005.600 5058.035 3020.400 5082.985 ;
      LAYER met5 ;
        RECT 3022.000 5058.035 3024.000 5082.985 ;
      LAYER met5 ;
        RECT 3025.600 5058.035 3040.400 5082.985 ;
      LAYER met5 ;
        RECT 3042.000 5058.035 3044.000 5082.985 ;
      LAYER met5 ;
        RECT 3045.600 5058.035 3060.400 5082.985 ;
      LAYER met5 ;
        RECT 3062.000 5058.035 3064.000 5082.985 ;
      LAYER met5 ;
        RECT 3065.600 5058.035 3080.400 5082.985 ;
      LAYER met5 ;
        RECT 3082.000 5058.035 3084.000 5082.985 ;
      LAYER met5 ;
        RECT 3085.600 5058.035 3100.400 5082.985 ;
      LAYER met5 ;
        RECT 3102.000 5058.035 3104.000 5082.985 ;
      LAYER met5 ;
        RECT 3105.600 5058.035 3120.400 5082.985 ;
      LAYER met5 ;
        RECT 3122.000 5058.035 3124.000 5082.985 ;
      LAYER met5 ;
        RECT 3125.600 5058.035 3140.400 5082.985 ;
      LAYER met5 ;
        RECT 3142.000 5058.035 3144.000 5082.985 ;
      LAYER met5 ;
        RECT 3145.600 5058.035 3160.400 5082.985 ;
      LAYER met5 ;
        RECT 3162.000 5058.035 3164.000 5082.985 ;
      LAYER met5 ;
        RECT 3165.600 5058.035 3180.400 5082.985 ;
      LAYER met5 ;
        RECT 3182.000 5058.035 3184.000 5082.985 ;
      LAYER met5 ;
        RECT 3185.600 5058.035 3200.400 5082.985 ;
      LAYER met5 ;
        RECT 3202.000 5058.035 3204.000 5082.985 ;
      LAYER met5 ;
        RECT 3205.600 5058.035 3220.400 5082.985 ;
      LAYER met5 ;
        RECT 3222.000 5058.035 3224.000 5082.985 ;
      LAYER met5 ;
        RECT 3225.600 5058.035 3240.400 5082.985 ;
      LAYER met5 ;
        RECT 3242.000 5058.035 3244.000 5082.985 ;
      LAYER met5 ;
        RECT 3245.600 5058.035 3260.400 5082.985 ;
      LAYER met5 ;
        RECT 3262.000 5058.035 3264.000 5082.985 ;
      LAYER met5 ;
        RECT 3265.600 5058.035 3280.400 5082.985 ;
      LAYER met5 ;
        RECT 3282.000 5058.035 3284.000 5082.985 ;
      LAYER met5 ;
        RECT 3285.600 5058.035 3300.400 5082.985 ;
      LAYER met5 ;
        RECT 3302.000 5058.035 3304.000 5082.985 ;
      LAYER met5 ;
        RECT 3305.600 5058.035 3320.400 5082.985 ;
      LAYER met5 ;
        RECT 3322.000 5058.035 3324.000 5082.985 ;
      LAYER met5 ;
        RECT 3325.600 5058.035 3340.400 5082.985 ;
      LAYER met5 ;
        RECT 3342.000 5058.035 3344.000 5082.985 ;
      LAYER met5 ;
        RECT 3345.600 5058.035 3360.400 5082.985 ;
      LAYER met5 ;
        RECT 3362.000 5058.035 3364.000 5082.985 ;
      LAYER met5 ;
        RECT 3365.600 5058.035 3380.400 5082.985 ;
      LAYER met5 ;
        RECT 3382.000 5058.035 3384.000 5082.985 ;
        RECT 3387.000 5058.035 3390.645 5082.985 ;
      LAYER met5 ;
        RECT 3392.245 5056.435 3588.000 5084.585 ;
      LAYER met5 ;
        RECT 2921.730 5052.185 3389.480 5056.435 ;
      LAYER met5 ;
        RECT 3391.080 5052.185 3588.000 5056.435 ;
      LAYER met5 ;
        RECT 2921.730 5046.335 3389.625 5050.585 ;
      LAYER met5 ;
        RECT 3391.225 5046.335 3588.000 5052.185 ;
      LAYER met5 ;
        RECT 2921.730 5035.735 3411.155 5044.735 ;
      LAYER met5 ;
        RECT 3412.755 5034.135 3588.000 5046.335 ;
      LAYER met5 ;
        RECT 2921.730 5029.685 3389.475 5034.135 ;
      LAYER met5 ;
        RECT 3391.075 5028.085 3588.000 5034.135 ;
      LAYER met5 ;
        RECT 2921.730 5024.840 3389.335 5028.085 ;
        RECT 2923.000 5024.835 3389.335 5024.840 ;
      LAYER met5 ;
        RECT 3390.935 5024.835 3588.000 5028.085 ;
      LAYER met5 ;
        RECT 2921.730 5019.985 3389.385 5023.235 ;
      LAYER met5 ;
        RECT 3390.985 5019.985 3588.000 5024.835 ;
      LAYER met5 ;
        RECT 2921.730 5013.935 3389.600 5018.385 ;
      LAYER met5 ;
        RECT 3391.200 5012.755 3588.000 5019.985 ;
        RECT 3391.200 5012.335 3434.135 5012.755 ;
      LAYER met5 ;
        RECT 2921.730 5007.885 3389.525 5012.335 ;
      LAYER met5 ;
        RECT 3391.125 5006.285 3434.135 5012.335 ;
        RECT 153.865 5003.035 201.145 5006.285 ;
      LAYER met5 ;
        RECT 202.745 5003.035 668.965 5006.285 ;
      LAYER met5 ;
        RECT 670.565 5003.035 745.370 5006.285 ;
      LAYER met5 ;
        RECT 746.970 5003.035 1213.965 5006.285 ;
      LAYER met5 ;
        RECT 1215.565 5003.035 1290.370 5006.285 ;
      LAYER met5 ;
        RECT 1291.970 5003.035 1758.965 5006.285 ;
      LAYER met5 ;
        RECT 1760.565 5003.035 1835.370 5006.285 ;
      LAYER met5 ;
        RECT 1836.970 5003.035 2303.965 5006.285 ;
      LAYER met5 ;
        RECT 2305.565 5003.035 2380.370 5006.285 ;
      LAYER met5 ;
        RECT 2381.970 5003.035 2848.965 5006.285 ;
      LAYER met5 ;
        RECT 2850.565 5003.035 2920.435 5006.285 ;
      LAYER met5 ;
        RECT 2922.035 5003.035 3389.470 5006.285 ;
      LAYER met5 ;
        RECT 3391.070 5003.035 3434.135 5006.285 ;
        RECT 153.865 4993.385 201.130 5003.035 ;
      LAYER met5 ;
        RECT 202.730 4996.985 669.270 5001.435 ;
      LAYER met5 ;
        RECT 153.865 4991.200 184.965 4993.385 ;
        RECT 192.615 4991.950 201.130 4993.385 ;
        RECT 153.865 4991.075 168.015 4991.200 ;
        RECT 175.665 4991.125 184.965 4991.200 ;
        RECT 159.915 4990.985 168.015 4991.075 ;
        RECT 181.715 4991.070 184.965 4991.125 ;
        RECT 159.915 4990.935 163.165 4990.985 ;
      LAYER met5 ;
        RECT 153.865 4457.730 158.315 4989.475 ;
        RECT 159.915 4459.000 163.165 4989.335 ;
        RECT 159.915 4457.730 163.160 4459.000 ;
        RECT 164.765 4457.730 168.015 4989.385 ;
        RECT 169.615 4457.730 174.065 4989.600 ;
        RECT 175.665 4457.730 180.115 4989.525 ;
        RECT 181.715 4458.035 184.965 4989.470 ;
        RECT 186.565 4457.730 191.015 4991.785 ;
        RECT 192.615 4457.730 197.865 4990.350 ;
      LAYER met5 ;
        RECT 199.465 4988.535 201.130 4991.950 ;
      LAYER met5 ;
        RECT 202.730 4990.135 669.270 4995.385 ;
      LAYER met5 ;
        RECT 670.870 4990.135 745.130 5003.035 ;
      LAYER met5 ;
        RECT 746.730 4996.985 1214.270 5001.435 ;
        RECT 746.730 4990.135 1214.270 4995.385 ;
      LAYER met5 ;
        RECT 1215.870 4990.135 1290.130 5003.035 ;
      LAYER met5 ;
        RECT 1291.730 4996.985 1759.270 5001.435 ;
        RECT 1291.730 4990.135 1759.270 4995.385 ;
      LAYER met5 ;
        RECT 1760.870 4990.135 1835.130 5003.035 ;
      LAYER met5 ;
        RECT 1836.730 4996.985 2304.270 5001.435 ;
        RECT 1836.730 4990.135 2304.270 4995.385 ;
      LAYER met5 ;
        RECT 2305.870 4990.135 2380.130 5003.035 ;
      LAYER met5 ;
        RECT 2381.730 4996.985 2849.270 5001.435 ;
        RECT 2381.730 4990.135 2849.270 4995.385 ;
      LAYER met5 ;
        RECT 2850.870 4990.135 2920.130 5003.035 ;
      LAYER met5 ;
        RECT 2921.730 4996.985 3391.785 5001.435 ;
      LAYER met5 ;
        RECT 3393.385 4995.385 3434.135 5003.035 ;
      LAYER met5 ;
        RECT 2921.730 4990.135 3390.350 4995.385 ;
      LAYER met5 ;
        RECT 3391.950 4988.535 3434.135 4995.385 ;
        RECT 199.465 4988.000 204.000 4988.535 ;
        RECT 3388.000 4986.870 3434.135 4988.535 ;
        RECT 3388.000 4984.000 3388.535 4986.870 ;
        RECT 3403.035 4986.855 3406.285 4986.870 ;
        RECT 181.715 4456.130 184.965 4456.435 ;
        RECT 0.000 4454.400 197.865 4456.130 ;
        RECT 0.000 4388.500 31.775 4454.400 ;
        RECT 97.590 4388.500 197.865 4454.400 ;
      LAYER met5 ;
        RECT 3390.135 4453.730 3395.385 4985.270 ;
        RECT 3396.985 4453.730 3401.435 4985.270 ;
        RECT 3403.035 4454.035 3406.285 4985.255 ;
        RECT 3407.885 4453.730 3412.335 4985.270 ;
        RECT 3413.935 4453.730 3418.385 4985.270 ;
        RECT 3419.985 4453.730 3423.235 4985.270 ;
        RECT 3424.840 4984.000 3428.085 4985.270 ;
        RECT 3424.835 4455.000 3428.085 4984.000 ;
        RECT 3424.840 4453.730 3428.085 4455.000 ;
        RECT 3429.685 4453.730 3434.135 4985.270 ;
        RECT 3435.735 4453.730 3444.735 5011.155 ;
      LAYER met5 ;
        RECT 3446.335 4987.455 3588.000 5012.755 ;
        RECT 3446.335 4986.870 3456.435 4987.455 ;
      LAYER met5 ;
        RECT 3446.335 4453.730 3450.585 4985.270 ;
        RECT 3452.185 4453.730 3456.435 4985.270 ;
        RECT 3458.035 4979.000 3482.985 4985.855 ;
      LAYER met5 ;
        RECT 3484.585 4984.000 3588.000 4987.455 ;
      LAYER met5 ;
        RECT 3458.035 4974.000 3482.985 4976.000 ;
      LAYER met5 ;
        RECT 3458.035 4957.600 3482.985 4972.400 ;
      LAYER met5 ;
        RECT 3458.035 4954.000 3482.985 4956.000 ;
      LAYER met5 ;
        RECT 3458.035 4937.600 3482.985 4952.400 ;
      LAYER met5 ;
        RECT 3458.035 4934.000 3482.985 4936.000 ;
      LAYER met5 ;
        RECT 3458.035 4917.600 3482.985 4932.400 ;
      LAYER met5 ;
        RECT 3458.035 4914.000 3482.985 4916.000 ;
      LAYER met5 ;
        RECT 3458.035 4897.600 3482.985 4912.400 ;
      LAYER met5 ;
        RECT 3458.035 4894.000 3482.985 4896.000 ;
      LAYER met5 ;
        RECT 3458.035 4877.600 3482.985 4892.400 ;
      LAYER met5 ;
        RECT 3458.035 4874.000 3482.985 4876.000 ;
      LAYER met5 ;
        RECT 3458.035 4857.600 3482.985 4872.400 ;
      LAYER met5 ;
        RECT 3458.035 4854.000 3482.985 4856.000 ;
      LAYER met5 ;
        RECT 3458.035 4837.600 3482.985 4852.400 ;
      LAYER met5 ;
        RECT 3458.035 4834.000 3482.985 4836.000 ;
      LAYER met5 ;
        RECT 3458.035 4817.600 3482.985 4832.400 ;
      LAYER met5 ;
        RECT 3458.035 4814.000 3482.985 4816.000 ;
      LAYER met5 ;
        RECT 3458.035 4797.600 3482.985 4812.400 ;
      LAYER met5 ;
        RECT 3458.035 4794.000 3482.985 4796.000 ;
      LAYER met5 ;
        RECT 3458.035 4777.600 3482.985 4792.400 ;
      LAYER met5 ;
        RECT 3458.035 4774.000 3482.985 4776.000 ;
      LAYER met5 ;
        RECT 3458.035 4757.600 3482.985 4772.400 ;
      LAYER met5 ;
        RECT 3458.035 4754.000 3482.985 4756.000 ;
      LAYER met5 ;
        RECT 3458.035 4737.600 3482.985 4752.400 ;
      LAYER met5 ;
        RECT 3458.035 4734.000 3482.985 4736.000 ;
      LAYER met5 ;
        RECT 3458.035 4717.600 3482.985 4732.400 ;
      LAYER met5 ;
        RECT 3458.035 4714.000 3482.985 4716.000 ;
      LAYER met5 ;
        RECT 3458.035 4697.600 3482.985 4712.400 ;
      LAYER met5 ;
        RECT 3458.035 4694.000 3482.985 4696.000 ;
      LAYER met5 ;
        RECT 3458.035 4677.600 3482.985 4692.400 ;
      LAYER met5 ;
        RECT 3458.035 4674.000 3482.985 4676.000 ;
      LAYER met5 ;
        RECT 3458.035 4657.600 3482.985 4672.400 ;
      LAYER met5 ;
        RECT 3458.035 4654.000 3482.985 4656.000 ;
      LAYER met5 ;
        RECT 3458.035 4637.600 3482.985 4652.400 ;
      LAYER met5 ;
        RECT 3458.035 4634.000 3482.985 4636.000 ;
      LAYER met5 ;
        RECT 3458.035 4617.600 3482.985 4632.400 ;
      LAYER met5 ;
        RECT 3458.035 4614.000 3482.985 4616.000 ;
      LAYER met5 ;
        RECT 3458.035 4597.600 3482.985 4612.400 ;
      LAYER met5 ;
        RECT 3458.035 4594.000 3482.985 4596.000 ;
      LAYER met5 ;
        RECT 3458.035 4577.600 3482.985 4592.400 ;
      LAYER met5 ;
        RECT 3458.035 4574.000 3482.985 4576.000 ;
      LAYER met5 ;
        RECT 3458.035 4557.600 3482.985 4572.400 ;
      LAYER met5 ;
        RECT 3458.035 4554.000 3482.985 4556.000 ;
      LAYER met5 ;
        RECT 3458.035 4537.600 3482.985 4552.400 ;
      LAYER met5 ;
        RECT 3458.035 4534.000 3482.985 4536.000 ;
      LAYER met5 ;
        RECT 3458.035 4517.600 3482.985 4532.400 ;
      LAYER met5 ;
        RECT 3458.035 4514.000 3482.985 4516.000 ;
      LAYER met5 ;
        RECT 3458.035 4497.600 3482.985 4512.400 ;
      LAYER met5 ;
        RECT 3458.035 4494.000 3482.985 4496.000 ;
      LAYER met5 ;
        RECT 3458.035 4477.600 3482.985 4492.400 ;
      LAYER met5 ;
        RECT 3458.035 4474.000 3482.985 4476.000 ;
      LAYER met5 ;
        RECT 3458.035 4457.600 3482.985 4472.400 ;
      LAYER met5 ;
        RECT 3458.035 4453.730 3482.985 4456.000 ;
        RECT 3563.785 4455.000 3588.000 4984.000 ;
      LAYER met5 ;
        RECT 3403.035 4452.130 3406.285 4452.435 ;
        RECT 3484.585 4452.130 3588.000 4455.000 ;
        RECT 0.000 4386.870 197.865 4388.500 ;
        RECT 3390.135 4447.285 3588.000 4452.130 ;
        RECT 3390.135 4387.445 3488.540 4447.285 ;
        RECT 3559.170 4387.445 3588.000 4447.285 ;
        RECT 0.000 4384.000 103.415 4386.870 ;
        RECT 181.715 4386.565 184.965 4386.870 ;
      LAYER met5 ;
        RECT 0.000 3855.000 24.215 4384.000 ;
        RECT 105.015 4379.000 129.965 4385.270 ;
        RECT 105.015 4374.000 129.965 4376.000 ;
      LAYER met5 ;
        RECT 105.015 4357.600 129.965 4372.400 ;
      LAYER met5 ;
        RECT 105.015 4354.000 129.965 4356.000 ;
      LAYER met5 ;
        RECT 105.015 4337.600 129.965 4352.400 ;
      LAYER met5 ;
        RECT 105.015 4334.000 129.965 4336.000 ;
      LAYER met5 ;
        RECT 105.015 4317.600 129.965 4332.400 ;
      LAYER met5 ;
        RECT 105.015 4314.000 129.965 4316.000 ;
      LAYER met5 ;
        RECT 105.015 4297.600 129.965 4312.400 ;
      LAYER met5 ;
        RECT 105.015 4294.000 129.965 4296.000 ;
      LAYER met5 ;
        RECT 105.015 4277.600 129.965 4292.400 ;
      LAYER met5 ;
        RECT 105.015 4274.000 129.965 4276.000 ;
      LAYER met5 ;
        RECT 105.015 4257.600 129.965 4272.400 ;
      LAYER met5 ;
        RECT 105.015 4254.000 129.965 4256.000 ;
      LAYER met5 ;
        RECT 105.015 4237.600 129.965 4252.400 ;
      LAYER met5 ;
        RECT 105.015 4234.000 129.965 4236.000 ;
      LAYER met5 ;
        RECT 105.015 4217.600 129.965 4232.400 ;
      LAYER met5 ;
        RECT 105.015 4214.000 129.965 4216.000 ;
      LAYER met5 ;
        RECT 105.015 4197.600 129.965 4212.400 ;
      LAYER met5 ;
        RECT 105.015 4194.000 129.965 4196.000 ;
      LAYER met5 ;
        RECT 105.015 4177.600 129.965 4192.400 ;
      LAYER met5 ;
        RECT 105.015 4174.000 129.965 4176.000 ;
      LAYER met5 ;
        RECT 105.015 4157.600 129.965 4172.400 ;
      LAYER met5 ;
        RECT 105.015 4154.000 129.965 4156.000 ;
      LAYER met5 ;
        RECT 105.015 4137.600 129.965 4152.400 ;
      LAYER met5 ;
        RECT 105.015 4134.000 129.965 4136.000 ;
      LAYER met5 ;
        RECT 105.015 4117.600 129.965 4132.400 ;
      LAYER met5 ;
        RECT 105.015 4114.000 129.965 4116.000 ;
      LAYER met5 ;
        RECT 105.015 4097.600 129.965 4112.400 ;
      LAYER met5 ;
        RECT 105.015 4094.000 129.965 4096.000 ;
      LAYER met5 ;
        RECT 105.015 4077.600 129.965 4092.400 ;
      LAYER met5 ;
        RECT 105.015 4074.000 129.965 4076.000 ;
      LAYER met5 ;
        RECT 105.015 4057.600 129.965 4072.400 ;
      LAYER met5 ;
        RECT 105.015 4054.000 129.965 4056.000 ;
      LAYER met5 ;
        RECT 105.015 4037.600 129.965 4052.400 ;
      LAYER met5 ;
        RECT 105.015 4034.000 129.965 4036.000 ;
      LAYER met5 ;
        RECT 105.015 4017.600 129.965 4032.400 ;
      LAYER met5 ;
        RECT 105.015 4014.000 129.965 4016.000 ;
      LAYER met5 ;
        RECT 105.015 3997.600 129.965 4012.400 ;
      LAYER met5 ;
        RECT 105.015 3994.000 129.965 3996.000 ;
      LAYER met5 ;
        RECT 105.015 3977.600 129.965 3992.400 ;
      LAYER met5 ;
        RECT 105.015 3974.000 129.965 3976.000 ;
      LAYER met5 ;
        RECT 105.015 3957.600 129.965 3972.400 ;
      LAYER met5 ;
        RECT 105.015 3954.000 129.965 3956.000 ;
      LAYER met5 ;
        RECT 105.015 3937.600 129.965 3952.400 ;
      LAYER met5 ;
        RECT 105.015 3934.000 129.965 3936.000 ;
      LAYER met5 ;
        RECT 105.015 3917.600 129.965 3932.400 ;
      LAYER met5 ;
        RECT 105.015 3914.000 129.965 3916.000 ;
      LAYER met5 ;
        RECT 105.015 3897.600 129.965 3912.400 ;
      LAYER met5 ;
        RECT 105.015 3894.000 129.965 3896.000 ;
      LAYER met5 ;
        RECT 105.015 3877.600 129.965 3892.400 ;
      LAYER met5 ;
        RECT 105.015 3874.000 129.965 3876.000 ;
      LAYER met5 ;
        RECT 105.015 3857.600 129.965 3872.400 ;
        RECT 0.000 3852.130 103.415 3855.000 ;
      LAYER met5 ;
        RECT 105.015 3853.730 129.965 3856.000 ;
        RECT 131.565 3853.730 135.815 4385.270 ;
        RECT 137.415 3853.730 141.665 4385.270 ;
        RECT 143.265 3853.730 152.265 4385.270 ;
        RECT 153.865 3853.730 158.315 4385.270 ;
        RECT 159.915 4384.000 163.160 4385.270 ;
        RECT 159.915 3855.000 163.165 4384.000 ;
        RECT 159.915 3853.730 163.160 3855.000 ;
        RECT 164.765 3853.730 168.015 4385.270 ;
        RECT 169.615 3853.730 174.065 4385.270 ;
        RECT 175.665 3853.730 180.115 4385.270 ;
        RECT 181.715 3853.970 184.965 4384.965 ;
        RECT 186.565 3853.730 191.015 4385.270 ;
        RECT 192.615 3853.730 197.865 4385.270 ;
      LAYER met5 ;
        RECT 3390.135 4382.870 3588.000 4387.445 ;
        RECT 3403.035 4382.565 3406.285 4382.870 ;
      LAYER met5 ;
        RECT 3380.660 4278.100 3383.180 4279.700 ;
        RECT 3380.660 4274.700 3382.260 4278.100 ;
      LAYER met5 ;
        RECT 181.715 3852.130 184.965 3852.370 ;
        RECT 0.000 3850.400 197.865 3852.130 ;
        RECT 0.000 3784.600 31.390 3850.400 ;
        RECT 97.040 3784.600 197.865 3850.400 ;
      LAYER met5 ;
        RECT 3390.135 3849.730 3395.385 4381.270 ;
        RECT 3396.985 3849.730 3401.435 4381.270 ;
        RECT 3403.035 3850.035 3406.285 4380.965 ;
        RECT 3407.885 3849.730 3412.335 4381.270 ;
        RECT 3413.935 3849.730 3418.385 4381.270 ;
        RECT 3419.985 3849.730 3423.235 4381.270 ;
        RECT 3424.840 4380.000 3428.085 4381.270 ;
        RECT 3424.835 3851.000 3428.085 4380.000 ;
        RECT 3424.840 3849.730 3428.085 3851.000 ;
        RECT 3429.685 3849.730 3434.135 4381.270 ;
        RECT 3435.735 3849.730 3444.735 4381.270 ;
        RECT 3446.335 3849.730 3450.585 4381.270 ;
        RECT 3452.185 3849.730 3456.435 4381.270 ;
        RECT 3458.035 4375.000 3482.985 4381.270 ;
      LAYER met5 ;
        RECT 3484.585 4380.000 3588.000 4382.870 ;
      LAYER met5 ;
        RECT 3458.035 4370.000 3482.985 4372.000 ;
      LAYER met5 ;
        RECT 3458.035 4353.600 3482.985 4368.400 ;
      LAYER met5 ;
        RECT 3458.035 4350.000 3482.985 4352.000 ;
      LAYER met5 ;
        RECT 3458.035 4333.600 3482.985 4348.400 ;
      LAYER met5 ;
        RECT 3458.035 4330.000 3482.985 4332.000 ;
      LAYER met5 ;
        RECT 3458.035 4313.600 3482.985 4328.400 ;
      LAYER met5 ;
        RECT 3458.035 4310.000 3482.985 4312.000 ;
      LAYER met5 ;
        RECT 3458.035 4293.600 3482.985 4308.400 ;
      LAYER met5 ;
        RECT 3458.035 4290.000 3482.985 4292.000 ;
      LAYER met5 ;
        RECT 3458.035 4273.600 3482.985 4288.400 ;
      LAYER met5 ;
        RECT 3458.035 4270.000 3482.985 4272.000 ;
      LAYER met5 ;
        RECT 3458.035 4253.600 3482.985 4268.400 ;
      LAYER met5 ;
        RECT 3458.035 4250.000 3482.985 4252.000 ;
      LAYER met5 ;
        RECT 3458.035 4233.600 3482.985 4248.400 ;
      LAYER met5 ;
        RECT 3458.035 4230.000 3482.985 4232.000 ;
      LAYER met5 ;
        RECT 3458.035 4213.600 3482.985 4228.400 ;
      LAYER met5 ;
        RECT 3458.035 4210.000 3482.985 4212.000 ;
      LAYER met5 ;
        RECT 3458.035 4193.600 3482.985 4208.400 ;
      LAYER met5 ;
        RECT 3458.035 4190.000 3482.985 4192.000 ;
      LAYER met5 ;
        RECT 3458.035 4173.600 3482.985 4188.400 ;
      LAYER met5 ;
        RECT 3458.035 4170.000 3482.985 4172.000 ;
      LAYER met5 ;
        RECT 3458.035 4153.600 3482.985 4168.400 ;
      LAYER met5 ;
        RECT 3458.035 4150.000 3482.985 4152.000 ;
      LAYER met5 ;
        RECT 3458.035 4133.600 3482.985 4148.400 ;
      LAYER met5 ;
        RECT 3458.035 4130.000 3482.985 4132.000 ;
      LAYER met5 ;
        RECT 3458.035 4113.600 3482.985 4128.400 ;
      LAYER met5 ;
        RECT 3458.035 4110.000 3482.985 4112.000 ;
      LAYER met5 ;
        RECT 3458.035 4093.600 3482.985 4108.400 ;
      LAYER met5 ;
        RECT 3458.035 4090.000 3482.985 4092.000 ;
      LAYER met5 ;
        RECT 3458.035 4073.600 3482.985 4088.400 ;
      LAYER met5 ;
        RECT 3458.035 4070.000 3482.985 4072.000 ;
      LAYER met5 ;
        RECT 3458.035 4053.600 3482.985 4068.400 ;
      LAYER met5 ;
        RECT 3458.035 4050.000 3482.985 4052.000 ;
      LAYER met5 ;
        RECT 3458.035 4033.600 3482.985 4048.400 ;
      LAYER met5 ;
        RECT 3458.035 4030.000 3482.985 4032.000 ;
      LAYER met5 ;
        RECT 3458.035 4013.600 3482.985 4028.400 ;
      LAYER met5 ;
        RECT 3458.035 4010.000 3482.985 4012.000 ;
      LAYER met5 ;
        RECT 3458.035 3993.600 3482.985 4008.400 ;
      LAYER met5 ;
        RECT 3458.035 3990.000 3482.985 3992.000 ;
      LAYER met5 ;
        RECT 3458.035 3973.600 3482.985 3988.400 ;
      LAYER met5 ;
        RECT 3458.035 3970.000 3482.985 3972.000 ;
      LAYER met5 ;
        RECT 3458.035 3953.600 3482.985 3968.400 ;
      LAYER met5 ;
        RECT 3458.035 3950.000 3482.985 3952.000 ;
      LAYER met5 ;
        RECT 3458.035 3933.600 3482.985 3948.400 ;
      LAYER met5 ;
        RECT 3458.035 3930.000 3482.985 3932.000 ;
      LAYER met5 ;
        RECT 3458.035 3913.600 3482.985 3928.400 ;
      LAYER met5 ;
        RECT 3458.035 3910.000 3482.985 3912.000 ;
      LAYER met5 ;
        RECT 3458.035 3893.600 3482.985 3908.400 ;
      LAYER met5 ;
        RECT 3458.035 3890.000 3482.985 3892.000 ;
      LAYER met5 ;
        RECT 3458.035 3873.600 3482.985 3888.400 ;
      LAYER met5 ;
        RECT 3458.035 3870.000 3482.985 3872.000 ;
      LAYER met5 ;
        RECT 3458.035 3853.600 3482.985 3868.400 ;
      LAYER met5 ;
        RECT 3458.035 3849.730 3482.985 3852.000 ;
        RECT 3563.785 3851.000 3588.000 4380.000 ;
      LAYER met5 ;
        RECT 3403.035 3848.130 3406.285 3848.435 ;
        RECT 3484.585 3848.130 3588.000 3851.000 ;
        RECT 3390.135 3841.400 3588.000 3848.130 ;
      LAYER met5 ;
        RECT 3380.660 3815.700 3387.780 3817.300 ;
      LAYER met5 ;
        RECT 0.000 3777.870 197.865 3784.600 ;
        RECT 0.000 3775.000 103.415 3777.870 ;
        RECT 181.715 3777.565 184.965 3777.870 ;
      LAYER met5 ;
        RECT 0.000 3247.000 24.215 3775.000 ;
        RECT 105.015 3771.000 129.965 3776.270 ;
        RECT 105.015 3766.000 129.965 3768.000 ;
      LAYER met5 ;
        RECT 105.015 3749.600 129.965 3764.400 ;
      LAYER met5 ;
        RECT 105.015 3746.000 129.965 3748.000 ;
      LAYER met5 ;
        RECT 105.015 3729.600 129.965 3744.400 ;
      LAYER met5 ;
        RECT 105.015 3726.000 129.965 3728.000 ;
      LAYER met5 ;
        RECT 105.015 3709.600 129.965 3724.400 ;
      LAYER met5 ;
        RECT 105.015 3706.000 129.965 3708.000 ;
      LAYER met5 ;
        RECT 105.015 3689.600 129.965 3704.400 ;
      LAYER met5 ;
        RECT 105.015 3686.000 129.965 3688.000 ;
      LAYER met5 ;
        RECT 105.015 3669.600 129.965 3684.400 ;
      LAYER met5 ;
        RECT 105.015 3666.000 129.965 3668.000 ;
      LAYER met5 ;
        RECT 105.015 3649.600 129.965 3664.400 ;
      LAYER met5 ;
        RECT 105.015 3646.000 129.965 3648.000 ;
      LAYER met5 ;
        RECT 105.015 3629.600 129.965 3644.400 ;
      LAYER met5 ;
        RECT 105.015 3626.000 129.965 3628.000 ;
      LAYER met5 ;
        RECT 105.015 3609.600 129.965 3624.400 ;
      LAYER met5 ;
        RECT 105.015 3606.000 129.965 3608.000 ;
      LAYER met5 ;
        RECT 105.015 3589.600 129.965 3604.400 ;
      LAYER met5 ;
        RECT 105.015 3586.000 129.965 3588.000 ;
      LAYER met5 ;
        RECT 105.015 3569.600 129.965 3584.400 ;
      LAYER met5 ;
        RECT 105.015 3566.000 129.965 3568.000 ;
      LAYER met5 ;
        RECT 105.015 3549.600 129.965 3564.400 ;
      LAYER met5 ;
        RECT 105.015 3546.000 129.965 3548.000 ;
      LAYER met5 ;
        RECT 105.015 3529.600 129.965 3544.400 ;
      LAYER met5 ;
        RECT 105.015 3526.000 129.965 3528.000 ;
      LAYER met5 ;
        RECT 105.015 3509.600 129.965 3524.400 ;
      LAYER met5 ;
        RECT 105.015 3506.000 129.965 3508.000 ;
      LAYER met5 ;
        RECT 105.015 3489.600 129.965 3504.400 ;
      LAYER met5 ;
        RECT 105.015 3486.000 129.965 3488.000 ;
      LAYER met5 ;
        RECT 105.015 3469.600 129.965 3484.400 ;
      LAYER met5 ;
        RECT 105.015 3466.000 129.965 3468.000 ;
      LAYER met5 ;
        RECT 105.015 3449.600 129.965 3464.400 ;
      LAYER met5 ;
        RECT 105.015 3446.000 129.965 3448.000 ;
      LAYER met5 ;
        RECT 105.015 3429.600 129.965 3444.400 ;
      LAYER met5 ;
        RECT 105.015 3426.000 129.965 3428.000 ;
      LAYER met5 ;
        RECT 105.015 3409.600 129.965 3424.400 ;
      LAYER met5 ;
        RECT 105.015 3406.000 129.965 3408.000 ;
      LAYER met5 ;
        RECT 105.015 3389.600 129.965 3404.400 ;
      LAYER met5 ;
        RECT 105.015 3386.000 129.965 3388.000 ;
      LAYER met5 ;
        RECT 105.015 3369.600 129.965 3384.400 ;
      LAYER met5 ;
        RECT 105.015 3366.000 129.965 3368.000 ;
      LAYER met5 ;
        RECT 105.015 3349.600 129.965 3364.400 ;
      LAYER met5 ;
        RECT 105.015 3346.000 129.965 3348.000 ;
      LAYER met5 ;
        RECT 105.015 3329.600 129.965 3344.400 ;
      LAYER met5 ;
        RECT 105.015 3326.000 129.965 3328.000 ;
      LAYER met5 ;
        RECT 105.015 3309.600 129.965 3324.400 ;
      LAYER met5 ;
        RECT 105.015 3306.000 129.965 3308.000 ;
      LAYER met5 ;
        RECT 105.015 3289.600 129.965 3304.400 ;
      LAYER met5 ;
        RECT 105.015 3286.000 129.965 3288.000 ;
      LAYER met5 ;
        RECT 105.015 3269.600 129.965 3284.400 ;
      LAYER met5 ;
        RECT 105.015 3266.000 129.965 3268.000 ;
      LAYER met5 ;
        RECT 105.015 3249.600 129.965 3264.400 ;
        RECT 0.000 3244.130 103.415 3247.000 ;
      LAYER met5 ;
        RECT 105.015 3245.730 129.965 3248.000 ;
        RECT 131.565 3245.730 135.815 3776.270 ;
        RECT 137.415 3245.730 141.665 3776.270 ;
        RECT 143.265 3245.730 152.265 3776.270 ;
        RECT 153.865 3245.730 158.315 3776.270 ;
        RECT 159.915 3775.000 163.160 3776.270 ;
        RECT 159.915 3247.000 163.165 3775.000 ;
        RECT 159.915 3245.730 163.160 3247.000 ;
        RECT 164.765 3245.730 168.015 3776.270 ;
        RECT 169.615 3245.730 174.065 3776.270 ;
        RECT 175.665 3245.730 180.115 3776.270 ;
        RECT 181.715 3245.970 184.965 3775.965 ;
        RECT 186.565 3245.730 191.015 3776.270 ;
        RECT 192.615 3245.730 197.865 3776.270 ;
      LAYER met5 ;
        RECT 3390.135 3775.600 3490.960 3841.400 ;
        RECT 3556.610 3775.600 3588.000 3841.400 ;
        RECT 3390.135 3773.870 3588.000 3775.600 ;
        RECT 3403.035 3773.630 3406.285 3773.870 ;
      LAYER met5 ;
        RECT 3382.500 3574.300 3386.860 3575.900 ;
      LAYER met5 ;
        RECT 181.715 3244.130 184.965 3244.370 ;
        RECT 0.000 3242.400 197.865 3244.130 ;
        RECT 0.000 3176.600 31.390 3242.400 ;
        RECT 97.040 3176.600 197.865 3242.400 ;
      LAYER met5 ;
        RECT 3390.135 3241.730 3395.385 3772.270 ;
        RECT 3396.985 3241.730 3401.435 3772.270 ;
        RECT 3403.035 3242.035 3406.285 3772.030 ;
        RECT 3407.885 3241.730 3412.335 3772.270 ;
        RECT 3413.935 3241.730 3418.385 3772.270 ;
        RECT 3419.985 3241.730 3423.235 3772.270 ;
        RECT 3424.840 3771.000 3428.085 3772.270 ;
        RECT 3424.835 3243.000 3428.085 3771.000 ;
        RECT 3424.840 3241.730 3428.085 3243.000 ;
        RECT 3429.685 3241.730 3434.135 3772.270 ;
        RECT 3435.735 3241.730 3444.735 3772.270 ;
        RECT 3446.335 3241.730 3450.585 3772.270 ;
        RECT 3452.185 3241.730 3456.435 3772.270 ;
        RECT 3458.035 3767.000 3482.985 3772.270 ;
      LAYER met5 ;
        RECT 3484.585 3771.000 3588.000 3773.870 ;
      LAYER met5 ;
        RECT 3458.035 3762.000 3482.985 3764.000 ;
      LAYER met5 ;
        RECT 3458.035 3745.600 3482.985 3760.400 ;
      LAYER met5 ;
        RECT 3458.035 3742.000 3482.985 3744.000 ;
      LAYER met5 ;
        RECT 3458.035 3725.600 3482.985 3740.400 ;
      LAYER met5 ;
        RECT 3458.035 3722.000 3482.985 3724.000 ;
      LAYER met5 ;
        RECT 3458.035 3705.600 3482.985 3720.400 ;
      LAYER met5 ;
        RECT 3458.035 3702.000 3482.985 3704.000 ;
      LAYER met5 ;
        RECT 3458.035 3685.600 3482.985 3700.400 ;
      LAYER met5 ;
        RECT 3458.035 3682.000 3482.985 3684.000 ;
      LAYER met5 ;
        RECT 3458.035 3665.600 3482.985 3680.400 ;
      LAYER met5 ;
        RECT 3458.035 3662.000 3482.985 3664.000 ;
      LAYER met5 ;
        RECT 3458.035 3645.600 3482.985 3660.400 ;
      LAYER met5 ;
        RECT 3458.035 3642.000 3482.985 3644.000 ;
      LAYER met5 ;
        RECT 3458.035 3625.600 3482.985 3640.400 ;
      LAYER met5 ;
        RECT 3458.035 3622.000 3482.985 3624.000 ;
      LAYER met5 ;
        RECT 3458.035 3605.600 3482.985 3620.400 ;
      LAYER met5 ;
        RECT 3458.035 3602.000 3482.985 3604.000 ;
      LAYER met5 ;
        RECT 3458.035 3585.600 3482.985 3600.400 ;
      LAYER met5 ;
        RECT 3458.035 3582.000 3482.985 3584.000 ;
      LAYER met5 ;
        RECT 3458.035 3565.600 3482.985 3580.400 ;
      LAYER met5 ;
        RECT 3458.035 3562.000 3482.985 3564.000 ;
      LAYER met5 ;
        RECT 3458.035 3545.600 3482.985 3560.400 ;
      LAYER met5 ;
        RECT 3458.035 3542.000 3482.985 3544.000 ;
      LAYER met5 ;
        RECT 3458.035 3525.600 3482.985 3540.400 ;
      LAYER met5 ;
        RECT 3458.035 3522.000 3482.985 3524.000 ;
      LAYER met5 ;
        RECT 3458.035 3505.600 3482.985 3520.400 ;
      LAYER met5 ;
        RECT 3458.035 3502.000 3482.985 3504.000 ;
      LAYER met5 ;
        RECT 3458.035 3485.600 3482.985 3500.400 ;
      LAYER met5 ;
        RECT 3458.035 3482.000 3482.985 3484.000 ;
      LAYER met5 ;
        RECT 3458.035 3465.600 3482.985 3480.400 ;
      LAYER met5 ;
        RECT 3458.035 3462.000 3482.985 3464.000 ;
      LAYER met5 ;
        RECT 3458.035 3445.600 3482.985 3460.400 ;
      LAYER met5 ;
        RECT 3458.035 3442.000 3482.985 3444.000 ;
      LAYER met5 ;
        RECT 3458.035 3425.600 3482.985 3440.400 ;
      LAYER met5 ;
        RECT 3458.035 3422.000 3482.985 3424.000 ;
      LAYER met5 ;
        RECT 3458.035 3405.600 3482.985 3420.400 ;
      LAYER met5 ;
        RECT 3458.035 3402.000 3482.985 3404.000 ;
      LAYER met5 ;
        RECT 3458.035 3385.600 3482.985 3400.400 ;
      LAYER met5 ;
        RECT 3458.035 3382.000 3482.985 3384.000 ;
      LAYER met5 ;
        RECT 3458.035 3365.600 3482.985 3380.400 ;
      LAYER met5 ;
        RECT 3458.035 3362.000 3482.985 3364.000 ;
      LAYER met5 ;
        RECT 3458.035 3345.600 3482.985 3360.400 ;
      LAYER met5 ;
        RECT 3458.035 3342.000 3482.985 3344.000 ;
      LAYER met5 ;
        RECT 3458.035 3325.600 3482.985 3340.400 ;
      LAYER met5 ;
        RECT 3458.035 3322.000 3482.985 3324.000 ;
      LAYER met5 ;
        RECT 3458.035 3305.600 3482.985 3320.400 ;
      LAYER met5 ;
        RECT 3458.035 3302.000 3482.985 3304.000 ;
      LAYER met5 ;
        RECT 3458.035 3285.600 3482.985 3300.400 ;
      LAYER met5 ;
        RECT 3458.035 3282.000 3482.985 3284.000 ;
      LAYER met5 ;
        RECT 3458.035 3265.600 3482.985 3280.400 ;
      LAYER met5 ;
        RECT 3458.035 3262.000 3482.985 3264.000 ;
      LAYER met5 ;
        RECT 3458.035 3245.600 3482.985 3260.400 ;
      LAYER met5 ;
        RECT 3458.035 3241.730 3482.985 3244.000 ;
        RECT 3563.785 3243.000 3588.000 3771.000 ;
      LAYER met5 ;
        RECT 3403.035 3240.130 3406.285 3240.435 ;
        RECT 3484.585 3240.130 3588.000 3243.000 ;
        RECT 0.000 3169.870 197.865 3176.600 ;
        RECT 3390.135 3233.400 3588.000 3240.130 ;
        RECT 0.000 3167.000 103.415 3169.870 ;
        RECT 181.715 3169.565 184.965 3169.870 ;
      LAYER met5 ;
        RECT 0.000 2638.000 24.215 3167.000 ;
        RECT 105.015 3162.000 129.965 3168.270 ;
        RECT 105.015 3157.000 129.965 3159.000 ;
      LAYER met5 ;
        RECT 105.015 3140.600 129.965 3155.400 ;
      LAYER met5 ;
        RECT 105.015 3137.000 129.965 3139.000 ;
      LAYER met5 ;
        RECT 105.015 3120.600 129.965 3135.400 ;
      LAYER met5 ;
        RECT 105.015 3117.000 129.965 3119.000 ;
      LAYER met5 ;
        RECT 105.015 3100.600 129.965 3115.400 ;
      LAYER met5 ;
        RECT 105.015 3097.000 129.965 3099.000 ;
      LAYER met5 ;
        RECT 105.015 3080.600 129.965 3095.400 ;
      LAYER met5 ;
        RECT 105.015 3077.000 129.965 3079.000 ;
      LAYER met5 ;
        RECT 105.015 3060.600 129.965 3075.400 ;
      LAYER met5 ;
        RECT 105.015 3057.000 129.965 3059.000 ;
      LAYER met5 ;
        RECT 105.015 3040.600 129.965 3055.400 ;
      LAYER met5 ;
        RECT 105.015 3037.000 129.965 3039.000 ;
      LAYER met5 ;
        RECT 105.015 3020.600 129.965 3035.400 ;
      LAYER met5 ;
        RECT 105.015 3017.000 129.965 3019.000 ;
      LAYER met5 ;
        RECT 105.015 3000.600 129.965 3015.400 ;
      LAYER met5 ;
        RECT 105.015 2997.000 129.965 2999.000 ;
      LAYER met5 ;
        RECT 105.015 2980.600 129.965 2995.400 ;
      LAYER met5 ;
        RECT 105.015 2977.000 129.965 2979.000 ;
      LAYER met5 ;
        RECT 105.015 2960.600 129.965 2975.400 ;
      LAYER met5 ;
        RECT 105.015 2957.000 129.965 2959.000 ;
      LAYER met5 ;
        RECT 105.015 2940.600 129.965 2955.400 ;
      LAYER met5 ;
        RECT 105.015 2937.000 129.965 2939.000 ;
      LAYER met5 ;
        RECT 105.015 2920.600 129.965 2935.400 ;
      LAYER met5 ;
        RECT 105.015 2917.000 129.965 2919.000 ;
      LAYER met5 ;
        RECT 105.015 2900.600 129.965 2915.400 ;
      LAYER met5 ;
        RECT 105.015 2897.000 129.965 2899.000 ;
      LAYER met5 ;
        RECT 105.015 2880.600 129.965 2895.400 ;
      LAYER met5 ;
        RECT 105.015 2877.000 129.965 2879.000 ;
      LAYER met5 ;
        RECT 105.015 2860.600 129.965 2875.400 ;
      LAYER met5 ;
        RECT 105.015 2857.000 129.965 2859.000 ;
      LAYER met5 ;
        RECT 105.015 2840.600 129.965 2855.400 ;
      LAYER met5 ;
        RECT 105.015 2837.000 129.965 2839.000 ;
      LAYER met5 ;
        RECT 105.015 2820.600 129.965 2835.400 ;
      LAYER met5 ;
        RECT 105.015 2817.000 129.965 2819.000 ;
      LAYER met5 ;
        RECT 105.015 2800.600 129.965 2815.400 ;
      LAYER met5 ;
        RECT 105.015 2797.000 129.965 2799.000 ;
      LAYER met5 ;
        RECT 105.015 2780.600 129.965 2795.400 ;
      LAYER met5 ;
        RECT 105.015 2777.000 129.965 2779.000 ;
      LAYER met5 ;
        RECT 105.015 2760.600 129.965 2775.400 ;
      LAYER met5 ;
        RECT 105.015 2757.000 129.965 2759.000 ;
      LAYER met5 ;
        RECT 105.015 2740.600 129.965 2755.400 ;
      LAYER met5 ;
        RECT 105.015 2737.000 129.965 2739.000 ;
      LAYER met5 ;
        RECT 105.015 2720.600 129.965 2735.400 ;
      LAYER met5 ;
        RECT 105.015 2717.000 129.965 2719.000 ;
      LAYER met5 ;
        RECT 105.015 2700.600 129.965 2715.400 ;
      LAYER met5 ;
        RECT 105.015 2697.000 129.965 2699.000 ;
      LAYER met5 ;
        RECT 105.015 2680.600 129.965 2695.400 ;
      LAYER met5 ;
        RECT 105.015 2677.000 129.965 2679.000 ;
      LAYER met5 ;
        RECT 105.015 2660.600 129.965 2675.400 ;
      LAYER met5 ;
        RECT 105.015 2657.000 129.965 2659.000 ;
      LAYER met5 ;
        RECT 105.015 2640.600 129.965 2655.400 ;
        RECT 0.000 2635.130 103.415 2638.000 ;
      LAYER met5 ;
        RECT 105.015 2636.730 129.965 2639.000 ;
        RECT 131.565 2636.730 135.815 3168.270 ;
        RECT 137.415 2636.730 141.665 3168.270 ;
        RECT 143.265 2636.730 152.265 3168.270 ;
        RECT 153.865 2636.730 158.315 3168.270 ;
        RECT 159.915 3167.000 163.160 3168.270 ;
        RECT 159.915 2638.000 163.165 3167.000 ;
        RECT 159.915 2636.730 163.160 2638.000 ;
        RECT 164.765 2636.730 168.015 3168.270 ;
        RECT 169.615 2636.730 174.065 3168.270 ;
        RECT 175.665 2636.730 180.115 3168.270 ;
        RECT 181.715 2636.970 184.965 3167.965 ;
        RECT 186.565 2636.730 191.015 3168.270 ;
        RECT 192.615 2636.730 197.865 3168.270 ;
      LAYER met5 ;
        RECT 3390.135 3167.600 3490.960 3233.400 ;
        RECT 3556.610 3167.600 3588.000 3233.400 ;
        RECT 3390.135 3165.870 3588.000 3167.600 ;
        RECT 3403.035 3165.630 3406.285 3165.870 ;
      LAYER met5 ;
        RECT 3380.660 2731.100 3387.780 2732.700 ;
        RECT 3380.660 2703.900 3386.860 2705.500 ;
      LAYER met5 ;
        RECT 181.715 2635.130 184.965 2635.370 ;
        RECT 0.000 2633.400 197.865 2635.130 ;
        RECT 0.000 2567.600 31.390 2633.400 ;
        RECT 97.040 2567.600 197.865 2633.400 ;
      LAYER met5 ;
        RECT 3390.135 2632.730 3395.385 3164.270 ;
        RECT 3396.985 2632.730 3401.435 3164.270 ;
        RECT 3403.035 2633.035 3406.285 3164.030 ;
        RECT 3407.885 2632.730 3412.335 3164.270 ;
        RECT 3413.935 2632.730 3418.385 3164.270 ;
        RECT 3419.985 2632.730 3423.235 3164.270 ;
        RECT 3424.840 3163.000 3428.085 3164.270 ;
        RECT 3424.835 2634.000 3428.085 3163.000 ;
        RECT 3424.840 2632.730 3428.085 2634.000 ;
        RECT 3429.685 2632.730 3434.135 3164.270 ;
        RECT 3435.735 2632.730 3444.735 3164.270 ;
        RECT 3446.335 2632.730 3450.585 3164.270 ;
        RECT 3452.185 2632.730 3456.435 3164.270 ;
        RECT 3458.035 3158.000 3482.985 3164.270 ;
      LAYER met5 ;
        RECT 3484.585 3163.000 3588.000 3165.870 ;
      LAYER met5 ;
        RECT 3458.035 3153.000 3482.985 3155.000 ;
      LAYER met5 ;
        RECT 3458.035 3136.600 3482.985 3151.400 ;
      LAYER met5 ;
        RECT 3458.035 3133.000 3482.985 3135.000 ;
      LAYER met5 ;
        RECT 3458.035 3116.600 3482.985 3131.400 ;
      LAYER met5 ;
        RECT 3458.035 3113.000 3482.985 3115.000 ;
      LAYER met5 ;
        RECT 3458.035 3096.600 3482.985 3111.400 ;
      LAYER met5 ;
        RECT 3458.035 3093.000 3482.985 3095.000 ;
      LAYER met5 ;
        RECT 3458.035 3076.600 3482.985 3091.400 ;
      LAYER met5 ;
        RECT 3458.035 3073.000 3482.985 3075.000 ;
      LAYER met5 ;
        RECT 3458.035 3056.600 3482.985 3071.400 ;
      LAYER met5 ;
        RECT 3458.035 3053.000 3482.985 3055.000 ;
      LAYER met5 ;
        RECT 3458.035 3036.600 3482.985 3051.400 ;
      LAYER met5 ;
        RECT 3458.035 3033.000 3482.985 3035.000 ;
      LAYER met5 ;
        RECT 3458.035 3016.600 3482.985 3031.400 ;
      LAYER met5 ;
        RECT 3458.035 3013.000 3482.985 3015.000 ;
      LAYER met5 ;
        RECT 3458.035 2996.600 3482.985 3011.400 ;
      LAYER met5 ;
        RECT 3458.035 2993.000 3482.985 2995.000 ;
      LAYER met5 ;
        RECT 3458.035 2976.600 3482.985 2991.400 ;
      LAYER met5 ;
        RECT 3458.035 2973.000 3482.985 2975.000 ;
      LAYER met5 ;
        RECT 3458.035 2956.600 3482.985 2971.400 ;
      LAYER met5 ;
        RECT 3458.035 2953.000 3482.985 2955.000 ;
      LAYER met5 ;
        RECT 3458.035 2936.600 3482.985 2951.400 ;
      LAYER met5 ;
        RECT 3458.035 2933.000 3482.985 2935.000 ;
      LAYER met5 ;
        RECT 3458.035 2916.600 3482.985 2931.400 ;
      LAYER met5 ;
        RECT 3458.035 2913.000 3482.985 2915.000 ;
      LAYER met5 ;
        RECT 3458.035 2896.600 3482.985 2911.400 ;
      LAYER met5 ;
        RECT 3458.035 2893.000 3482.985 2895.000 ;
      LAYER met5 ;
        RECT 3458.035 2876.600 3482.985 2891.400 ;
      LAYER met5 ;
        RECT 3458.035 2873.000 3482.985 2875.000 ;
      LAYER met5 ;
        RECT 3458.035 2856.600 3482.985 2871.400 ;
      LAYER met5 ;
        RECT 3458.035 2853.000 3482.985 2855.000 ;
      LAYER met5 ;
        RECT 3458.035 2836.600 3482.985 2851.400 ;
      LAYER met5 ;
        RECT 3458.035 2833.000 3482.985 2835.000 ;
      LAYER met5 ;
        RECT 3458.035 2816.600 3482.985 2831.400 ;
      LAYER met5 ;
        RECT 3458.035 2813.000 3482.985 2815.000 ;
      LAYER met5 ;
        RECT 3458.035 2796.600 3482.985 2811.400 ;
      LAYER met5 ;
        RECT 3458.035 2793.000 3482.985 2795.000 ;
      LAYER met5 ;
        RECT 3458.035 2776.600 3482.985 2791.400 ;
      LAYER met5 ;
        RECT 3458.035 2773.000 3482.985 2775.000 ;
      LAYER met5 ;
        RECT 3458.035 2756.600 3482.985 2771.400 ;
      LAYER met5 ;
        RECT 3458.035 2753.000 3482.985 2755.000 ;
      LAYER met5 ;
        RECT 3458.035 2736.600 3482.985 2751.400 ;
      LAYER met5 ;
        RECT 3458.035 2733.000 3482.985 2735.000 ;
      LAYER met5 ;
        RECT 3458.035 2716.600 3482.985 2731.400 ;
      LAYER met5 ;
        RECT 3458.035 2713.000 3482.985 2715.000 ;
      LAYER met5 ;
        RECT 3458.035 2696.600 3482.985 2711.400 ;
      LAYER met5 ;
        RECT 3458.035 2693.000 3482.985 2695.000 ;
      LAYER met5 ;
        RECT 3458.035 2676.600 3482.985 2691.400 ;
      LAYER met5 ;
        RECT 3458.035 2673.000 3482.985 2675.000 ;
      LAYER met5 ;
        RECT 3458.035 2656.600 3482.985 2671.400 ;
      LAYER met5 ;
        RECT 3458.035 2653.000 3482.985 2655.000 ;
      LAYER met5 ;
        RECT 3458.035 2636.600 3482.985 2651.400 ;
      LAYER met5 ;
        RECT 3458.035 2632.730 3482.985 2635.000 ;
        RECT 3563.785 2634.000 3588.000 3163.000 ;
      LAYER met5 ;
        RECT 3403.035 2631.130 3406.285 2631.435 ;
        RECT 3484.585 2631.130 3588.000 2634.000 ;
        RECT 0.000 2560.870 197.865 2567.600 ;
        RECT 3390.135 2624.400 3588.000 2631.130 ;
        RECT 0.000 2558.000 103.415 2560.870 ;
        RECT 181.715 2560.565 184.965 2560.870 ;
      LAYER met5 ;
        RECT 0.000 2029.000 24.215 2558.000 ;
        RECT 105.015 2553.000 129.965 2559.270 ;
        RECT 105.015 2548.000 129.965 2550.000 ;
      LAYER met5 ;
        RECT 105.015 2531.600 129.965 2546.400 ;
      LAYER met5 ;
        RECT 105.015 2528.000 129.965 2530.000 ;
      LAYER met5 ;
        RECT 105.015 2511.600 129.965 2526.400 ;
      LAYER met5 ;
        RECT 105.015 2508.000 129.965 2510.000 ;
      LAYER met5 ;
        RECT 105.015 2491.600 129.965 2506.400 ;
      LAYER met5 ;
        RECT 105.015 2488.000 129.965 2490.000 ;
      LAYER met5 ;
        RECT 105.015 2471.600 129.965 2486.400 ;
      LAYER met5 ;
        RECT 105.015 2468.000 129.965 2470.000 ;
      LAYER met5 ;
        RECT 105.015 2451.600 129.965 2466.400 ;
      LAYER met5 ;
        RECT 105.015 2448.000 129.965 2450.000 ;
      LAYER met5 ;
        RECT 105.015 2431.600 129.965 2446.400 ;
      LAYER met5 ;
        RECT 105.015 2428.000 129.965 2430.000 ;
      LAYER met5 ;
        RECT 105.015 2411.600 129.965 2426.400 ;
      LAYER met5 ;
        RECT 105.015 2408.000 129.965 2410.000 ;
      LAYER met5 ;
        RECT 105.015 2391.600 129.965 2406.400 ;
      LAYER met5 ;
        RECT 105.015 2388.000 129.965 2390.000 ;
      LAYER met5 ;
        RECT 105.015 2371.600 129.965 2386.400 ;
      LAYER met5 ;
        RECT 105.015 2368.000 129.965 2370.000 ;
      LAYER met5 ;
        RECT 105.015 2351.600 129.965 2366.400 ;
      LAYER met5 ;
        RECT 105.015 2348.000 129.965 2350.000 ;
      LAYER met5 ;
        RECT 105.015 2331.600 129.965 2346.400 ;
      LAYER met5 ;
        RECT 105.015 2328.000 129.965 2330.000 ;
      LAYER met5 ;
        RECT 105.015 2311.600 129.965 2326.400 ;
      LAYER met5 ;
        RECT 105.015 2308.000 129.965 2310.000 ;
      LAYER met5 ;
        RECT 105.015 2291.600 129.965 2306.400 ;
      LAYER met5 ;
        RECT 105.015 2288.000 129.965 2290.000 ;
      LAYER met5 ;
        RECT 105.015 2271.600 129.965 2286.400 ;
      LAYER met5 ;
        RECT 105.015 2268.000 129.965 2270.000 ;
      LAYER met5 ;
        RECT 105.015 2251.600 129.965 2266.400 ;
      LAYER met5 ;
        RECT 105.015 2248.000 129.965 2250.000 ;
      LAYER met5 ;
        RECT 105.015 2231.600 129.965 2246.400 ;
      LAYER met5 ;
        RECT 105.015 2228.000 129.965 2230.000 ;
      LAYER met5 ;
        RECT 105.015 2211.600 129.965 2226.400 ;
      LAYER met5 ;
        RECT 105.015 2208.000 129.965 2210.000 ;
      LAYER met5 ;
        RECT 105.015 2191.600 129.965 2206.400 ;
      LAYER met5 ;
        RECT 105.015 2188.000 129.965 2190.000 ;
      LAYER met5 ;
        RECT 105.015 2171.600 129.965 2186.400 ;
      LAYER met5 ;
        RECT 105.015 2168.000 129.965 2170.000 ;
      LAYER met5 ;
        RECT 105.015 2151.600 129.965 2166.400 ;
      LAYER met5 ;
        RECT 105.015 2148.000 129.965 2150.000 ;
      LAYER met5 ;
        RECT 105.015 2131.600 129.965 2146.400 ;
      LAYER met5 ;
        RECT 105.015 2128.000 129.965 2130.000 ;
      LAYER met5 ;
        RECT 105.015 2111.600 129.965 2126.400 ;
      LAYER met5 ;
        RECT 105.015 2108.000 129.965 2110.000 ;
      LAYER met5 ;
        RECT 105.015 2091.600 129.965 2106.400 ;
      LAYER met5 ;
        RECT 105.015 2088.000 129.965 2090.000 ;
      LAYER met5 ;
        RECT 105.015 2071.600 129.965 2086.400 ;
      LAYER met5 ;
        RECT 105.015 2068.000 129.965 2070.000 ;
      LAYER met5 ;
        RECT 105.015 2051.600 129.965 2066.400 ;
      LAYER met5 ;
        RECT 105.015 2048.000 129.965 2050.000 ;
      LAYER met5 ;
        RECT 105.015 2031.600 129.965 2046.400 ;
        RECT 0.000 2026.130 103.415 2029.000 ;
      LAYER met5 ;
        RECT 105.015 2027.730 129.965 2030.000 ;
        RECT 131.565 2027.730 135.815 2559.270 ;
        RECT 137.415 2027.730 141.665 2559.270 ;
        RECT 143.265 2027.730 152.265 2559.270 ;
        RECT 153.865 2027.730 158.315 2559.270 ;
        RECT 159.915 2558.000 163.160 2559.270 ;
        RECT 159.915 2029.000 163.165 2558.000 ;
        RECT 159.915 2027.730 163.160 2029.000 ;
        RECT 164.765 2027.730 168.015 2559.270 ;
        RECT 169.615 2027.730 174.065 2559.270 ;
        RECT 175.665 2027.730 180.115 2559.270 ;
        RECT 181.715 2027.970 184.965 2558.965 ;
        RECT 186.565 2027.730 191.015 2559.270 ;
        RECT 192.615 2027.730 197.865 2559.270 ;
      LAYER met5 ;
        RECT 3390.135 2558.600 3490.960 2624.400 ;
        RECT 3556.610 2558.600 3588.000 2624.400 ;
        RECT 3390.135 2556.870 3588.000 2558.600 ;
        RECT 3403.035 2556.630 3406.285 2556.870 ;
        RECT 181.715 2026.130 184.965 2026.370 ;
        RECT 0.000 2024.400 197.865 2026.130 ;
        RECT 0.000 1958.600 31.390 2024.400 ;
        RECT 97.040 1958.600 197.865 2024.400 ;
      LAYER met5 ;
        RECT 3390.135 2023.730 3395.385 2555.270 ;
        RECT 3396.985 2023.730 3401.435 2555.270 ;
        RECT 3403.035 2024.035 3406.285 2555.030 ;
        RECT 3407.885 2023.730 3412.335 2555.270 ;
        RECT 3413.935 2023.730 3418.385 2555.270 ;
        RECT 3419.985 2023.730 3423.235 2555.270 ;
        RECT 3424.840 2554.000 3428.085 2555.270 ;
        RECT 3424.835 2025.000 3428.085 2554.000 ;
        RECT 3424.840 2023.730 3428.085 2025.000 ;
        RECT 3429.685 2023.730 3434.135 2555.270 ;
        RECT 3435.735 2023.730 3444.735 2555.270 ;
        RECT 3446.335 2023.730 3450.585 2555.270 ;
        RECT 3452.185 2023.730 3456.435 2555.270 ;
        RECT 3458.035 2549.000 3482.985 2555.270 ;
      LAYER met5 ;
        RECT 3484.585 2554.000 3588.000 2556.870 ;
      LAYER met5 ;
        RECT 3458.035 2544.000 3482.985 2546.000 ;
      LAYER met5 ;
        RECT 3458.035 2527.600 3482.985 2542.400 ;
      LAYER met5 ;
        RECT 3458.035 2524.000 3482.985 2526.000 ;
      LAYER met5 ;
        RECT 3458.035 2507.600 3482.985 2522.400 ;
      LAYER met5 ;
        RECT 3458.035 2504.000 3482.985 2506.000 ;
      LAYER met5 ;
        RECT 3458.035 2487.600 3482.985 2502.400 ;
      LAYER met5 ;
        RECT 3458.035 2484.000 3482.985 2486.000 ;
      LAYER met5 ;
        RECT 3458.035 2467.600 3482.985 2482.400 ;
      LAYER met5 ;
        RECT 3458.035 2464.000 3482.985 2466.000 ;
      LAYER met5 ;
        RECT 3458.035 2447.600 3482.985 2462.400 ;
      LAYER met5 ;
        RECT 3458.035 2444.000 3482.985 2446.000 ;
      LAYER met5 ;
        RECT 3458.035 2427.600 3482.985 2442.400 ;
      LAYER met5 ;
        RECT 3458.035 2424.000 3482.985 2426.000 ;
      LAYER met5 ;
        RECT 3458.035 2407.600 3482.985 2422.400 ;
      LAYER met5 ;
        RECT 3458.035 2404.000 3482.985 2406.000 ;
      LAYER met5 ;
        RECT 3458.035 2387.600 3482.985 2402.400 ;
      LAYER met5 ;
        RECT 3458.035 2384.000 3482.985 2386.000 ;
      LAYER met5 ;
        RECT 3458.035 2367.600 3482.985 2382.400 ;
      LAYER met5 ;
        RECT 3458.035 2364.000 3482.985 2366.000 ;
      LAYER met5 ;
        RECT 3458.035 2347.600 3482.985 2362.400 ;
      LAYER met5 ;
        RECT 3458.035 2344.000 3482.985 2346.000 ;
      LAYER met5 ;
        RECT 3458.035 2327.600 3482.985 2342.400 ;
      LAYER met5 ;
        RECT 3458.035 2324.000 3482.985 2326.000 ;
      LAYER met5 ;
        RECT 3458.035 2307.600 3482.985 2322.400 ;
      LAYER met5 ;
        RECT 3458.035 2304.000 3482.985 2306.000 ;
      LAYER met5 ;
        RECT 3458.035 2287.600 3482.985 2302.400 ;
      LAYER met5 ;
        RECT 3458.035 2284.000 3482.985 2286.000 ;
      LAYER met5 ;
        RECT 3458.035 2267.600 3482.985 2282.400 ;
      LAYER met5 ;
        RECT 3458.035 2264.000 3482.985 2266.000 ;
      LAYER met5 ;
        RECT 3458.035 2247.600 3482.985 2262.400 ;
      LAYER met5 ;
        RECT 3458.035 2244.000 3482.985 2246.000 ;
      LAYER met5 ;
        RECT 3458.035 2227.600 3482.985 2242.400 ;
      LAYER met5 ;
        RECT 3458.035 2224.000 3482.985 2226.000 ;
      LAYER met5 ;
        RECT 3458.035 2207.600 3482.985 2222.400 ;
      LAYER met5 ;
        RECT 3458.035 2204.000 3482.985 2206.000 ;
      LAYER met5 ;
        RECT 3458.035 2187.600 3482.985 2202.400 ;
      LAYER met5 ;
        RECT 3458.035 2184.000 3482.985 2186.000 ;
      LAYER met5 ;
        RECT 3458.035 2167.600 3482.985 2182.400 ;
      LAYER met5 ;
        RECT 3458.035 2164.000 3482.985 2166.000 ;
      LAYER met5 ;
        RECT 3458.035 2147.600 3482.985 2162.400 ;
      LAYER met5 ;
        RECT 3458.035 2144.000 3482.985 2146.000 ;
      LAYER met5 ;
        RECT 3458.035 2127.600 3482.985 2142.400 ;
      LAYER met5 ;
        RECT 3458.035 2124.000 3482.985 2126.000 ;
      LAYER met5 ;
        RECT 3458.035 2107.600 3482.985 2122.400 ;
      LAYER met5 ;
        RECT 3458.035 2104.000 3482.985 2106.000 ;
      LAYER met5 ;
        RECT 3458.035 2087.600 3482.985 2102.400 ;
      LAYER met5 ;
        RECT 3458.035 2084.000 3482.985 2086.000 ;
      LAYER met5 ;
        RECT 3458.035 2067.600 3482.985 2082.400 ;
      LAYER met5 ;
        RECT 3458.035 2064.000 3482.985 2066.000 ;
      LAYER met5 ;
        RECT 3458.035 2047.600 3482.985 2062.400 ;
      LAYER met5 ;
        RECT 3458.035 2044.000 3482.985 2046.000 ;
      LAYER met5 ;
        RECT 3458.035 2027.600 3482.985 2042.400 ;
      LAYER met5 ;
        RECT 3458.035 2023.730 3482.985 2026.000 ;
        RECT 3563.785 2025.000 3588.000 2554.000 ;
      LAYER met5 ;
        RECT 3403.035 2022.130 3406.285 2022.435 ;
        RECT 3484.585 2022.130 3588.000 2025.000 ;
        RECT 0.000 1951.870 197.865 1958.600 ;
        RECT 3390.135 2015.400 3588.000 2022.130 ;
        RECT 0.000 1949.000 103.415 1951.870 ;
        RECT 181.715 1951.565 184.965 1951.870 ;
      LAYER met5 ;
        RECT 0.000 1421.000 24.215 1949.000 ;
        RECT 105.015 1945.000 129.965 1950.270 ;
        RECT 105.015 1940.000 129.965 1942.000 ;
      LAYER met5 ;
        RECT 105.015 1923.600 129.965 1938.400 ;
      LAYER met5 ;
        RECT 105.015 1920.000 129.965 1922.000 ;
      LAYER met5 ;
        RECT 105.015 1903.600 129.965 1918.400 ;
      LAYER met5 ;
        RECT 105.015 1900.000 129.965 1902.000 ;
      LAYER met5 ;
        RECT 105.015 1883.600 129.965 1898.400 ;
      LAYER met5 ;
        RECT 105.015 1880.000 129.965 1882.000 ;
      LAYER met5 ;
        RECT 105.015 1863.600 129.965 1878.400 ;
      LAYER met5 ;
        RECT 105.015 1860.000 129.965 1862.000 ;
      LAYER met5 ;
        RECT 105.015 1843.600 129.965 1858.400 ;
      LAYER met5 ;
        RECT 105.015 1840.000 129.965 1842.000 ;
      LAYER met5 ;
        RECT 105.015 1823.600 129.965 1838.400 ;
      LAYER met5 ;
        RECT 105.015 1820.000 129.965 1822.000 ;
      LAYER met5 ;
        RECT 105.015 1803.600 129.965 1818.400 ;
      LAYER met5 ;
        RECT 105.015 1800.000 129.965 1802.000 ;
      LAYER met5 ;
        RECT 105.015 1783.600 129.965 1798.400 ;
      LAYER met5 ;
        RECT 105.015 1780.000 129.965 1782.000 ;
      LAYER met5 ;
        RECT 105.015 1763.600 129.965 1778.400 ;
      LAYER met5 ;
        RECT 105.015 1760.000 129.965 1762.000 ;
      LAYER met5 ;
        RECT 105.015 1743.600 129.965 1758.400 ;
      LAYER met5 ;
        RECT 105.015 1740.000 129.965 1742.000 ;
      LAYER met5 ;
        RECT 105.015 1723.600 129.965 1738.400 ;
      LAYER met5 ;
        RECT 105.015 1720.000 129.965 1722.000 ;
      LAYER met5 ;
        RECT 105.015 1703.600 129.965 1718.400 ;
      LAYER met5 ;
        RECT 105.015 1700.000 129.965 1702.000 ;
      LAYER met5 ;
        RECT 105.015 1683.600 129.965 1698.400 ;
      LAYER met5 ;
        RECT 105.015 1680.000 129.965 1682.000 ;
      LAYER met5 ;
        RECT 105.015 1663.600 129.965 1678.400 ;
      LAYER met5 ;
        RECT 105.015 1660.000 129.965 1662.000 ;
      LAYER met5 ;
        RECT 105.015 1643.600 129.965 1658.400 ;
      LAYER met5 ;
        RECT 105.015 1640.000 129.965 1642.000 ;
      LAYER met5 ;
        RECT 105.015 1623.600 129.965 1638.400 ;
      LAYER met5 ;
        RECT 105.015 1620.000 129.965 1622.000 ;
      LAYER met5 ;
        RECT 105.015 1603.600 129.965 1618.400 ;
      LAYER met5 ;
        RECT 105.015 1600.000 129.965 1602.000 ;
      LAYER met5 ;
        RECT 105.015 1583.600 129.965 1598.400 ;
      LAYER met5 ;
        RECT 105.015 1580.000 129.965 1582.000 ;
      LAYER met5 ;
        RECT 105.015 1563.600 129.965 1578.400 ;
      LAYER met5 ;
        RECT 105.015 1560.000 129.965 1562.000 ;
      LAYER met5 ;
        RECT 105.015 1543.600 129.965 1558.400 ;
      LAYER met5 ;
        RECT 105.015 1540.000 129.965 1542.000 ;
      LAYER met5 ;
        RECT 105.015 1523.600 129.965 1538.400 ;
      LAYER met5 ;
        RECT 105.015 1520.000 129.965 1522.000 ;
      LAYER met5 ;
        RECT 105.015 1503.600 129.965 1518.400 ;
      LAYER met5 ;
        RECT 105.015 1500.000 129.965 1502.000 ;
      LAYER met5 ;
        RECT 105.015 1483.600 129.965 1498.400 ;
      LAYER met5 ;
        RECT 105.015 1480.000 129.965 1482.000 ;
      LAYER met5 ;
        RECT 105.015 1463.600 129.965 1478.400 ;
      LAYER met5 ;
        RECT 105.015 1460.000 129.965 1462.000 ;
      LAYER met5 ;
        RECT 105.015 1443.600 129.965 1458.400 ;
      LAYER met5 ;
        RECT 105.015 1440.000 129.965 1442.000 ;
      LAYER met5 ;
        RECT 105.015 1423.600 129.965 1438.400 ;
        RECT 0.000 1418.130 103.415 1421.000 ;
      LAYER met5 ;
        RECT 105.015 1419.730 129.965 1422.000 ;
        RECT 131.565 1419.730 135.815 1950.270 ;
        RECT 137.415 1419.730 141.665 1950.270 ;
        RECT 143.265 1419.730 152.265 1950.270 ;
        RECT 153.865 1419.730 158.315 1950.270 ;
        RECT 159.915 1949.000 163.160 1950.270 ;
        RECT 159.915 1421.000 163.165 1949.000 ;
        RECT 159.915 1419.730 163.160 1421.000 ;
        RECT 164.765 1419.730 168.015 1950.270 ;
        RECT 169.615 1419.730 174.065 1950.270 ;
        RECT 175.665 1419.730 180.115 1950.270 ;
        RECT 181.715 1419.970 184.965 1949.965 ;
        RECT 186.565 1419.730 191.015 1950.270 ;
        RECT 192.615 1419.730 197.865 1950.270 ;
      LAYER met5 ;
        RECT 3390.135 1949.600 3490.960 2015.400 ;
        RECT 3556.610 1949.600 3588.000 2015.400 ;
        RECT 3390.135 1947.870 3588.000 1949.600 ;
        RECT 3403.035 1947.630 3406.285 1947.870 ;
      LAYER met5 ;
        RECT 3380.660 1864.100 3383.180 1865.700 ;
        RECT 3380.660 1860.700 3382.260 1864.100 ;
      LAYER met5 ;
        RECT 181.715 1418.130 184.965 1418.370 ;
        RECT 0.000 1416.400 197.865 1418.130 ;
        RECT 0.000 1350.600 31.390 1416.400 ;
        RECT 97.040 1350.600 197.865 1416.400 ;
      LAYER met5 ;
        RECT 3390.135 1415.730 3395.385 1946.270 ;
        RECT 3396.985 1415.730 3401.435 1946.270 ;
        RECT 3403.035 1416.035 3406.285 1946.030 ;
        RECT 3407.885 1415.730 3412.335 1946.270 ;
        RECT 3413.935 1415.730 3418.385 1946.270 ;
        RECT 3419.985 1415.730 3423.235 1946.270 ;
        RECT 3424.840 1945.000 3428.085 1946.270 ;
        RECT 3424.835 1417.000 3428.085 1945.000 ;
        RECT 3424.840 1415.730 3428.085 1417.000 ;
        RECT 3429.685 1415.730 3434.135 1946.270 ;
        RECT 3435.735 1415.730 3444.735 1946.270 ;
        RECT 3446.335 1415.730 3450.585 1946.270 ;
        RECT 3452.185 1415.730 3456.435 1946.270 ;
        RECT 3458.035 1941.000 3482.985 1946.270 ;
      LAYER met5 ;
        RECT 3484.585 1945.000 3588.000 1947.870 ;
      LAYER met5 ;
        RECT 3458.035 1936.000 3482.985 1938.000 ;
      LAYER met5 ;
        RECT 3458.035 1919.600 3482.985 1934.400 ;
      LAYER met5 ;
        RECT 3458.035 1916.000 3482.985 1918.000 ;
      LAYER met5 ;
        RECT 3458.035 1899.600 3482.985 1914.400 ;
      LAYER met5 ;
        RECT 3458.035 1896.000 3482.985 1898.000 ;
      LAYER met5 ;
        RECT 3458.035 1879.600 3482.985 1894.400 ;
      LAYER met5 ;
        RECT 3458.035 1876.000 3482.985 1878.000 ;
      LAYER met5 ;
        RECT 3458.035 1859.600 3482.985 1874.400 ;
      LAYER met5 ;
        RECT 3458.035 1856.000 3482.985 1858.000 ;
      LAYER met5 ;
        RECT 3458.035 1839.600 3482.985 1854.400 ;
      LAYER met5 ;
        RECT 3458.035 1836.000 3482.985 1838.000 ;
      LAYER met5 ;
        RECT 3458.035 1819.600 3482.985 1834.400 ;
      LAYER met5 ;
        RECT 3458.035 1816.000 3482.985 1818.000 ;
      LAYER met5 ;
        RECT 3458.035 1799.600 3482.985 1814.400 ;
      LAYER met5 ;
        RECT 3458.035 1796.000 3482.985 1798.000 ;
      LAYER met5 ;
        RECT 3458.035 1779.600 3482.985 1794.400 ;
      LAYER met5 ;
        RECT 3458.035 1776.000 3482.985 1778.000 ;
      LAYER met5 ;
        RECT 3458.035 1759.600 3482.985 1774.400 ;
      LAYER met5 ;
        RECT 3458.035 1756.000 3482.985 1758.000 ;
      LAYER met5 ;
        RECT 3458.035 1739.600 3482.985 1754.400 ;
      LAYER met5 ;
        RECT 3458.035 1736.000 3482.985 1738.000 ;
      LAYER met5 ;
        RECT 3458.035 1719.600 3482.985 1734.400 ;
      LAYER met5 ;
        RECT 3458.035 1716.000 3482.985 1718.000 ;
      LAYER met5 ;
        RECT 3458.035 1699.600 3482.985 1714.400 ;
      LAYER met5 ;
        RECT 3458.035 1696.000 3482.985 1698.000 ;
      LAYER met5 ;
        RECT 3458.035 1679.600 3482.985 1694.400 ;
      LAYER met5 ;
        RECT 3458.035 1676.000 3482.985 1678.000 ;
      LAYER met5 ;
        RECT 3458.035 1659.600 3482.985 1674.400 ;
      LAYER met5 ;
        RECT 3458.035 1656.000 3482.985 1658.000 ;
      LAYER met5 ;
        RECT 3458.035 1639.600 3482.985 1654.400 ;
      LAYER met5 ;
        RECT 3458.035 1636.000 3482.985 1638.000 ;
      LAYER met5 ;
        RECT 3458.035 1619.600 3482.985 1634.400 ;
      LAYER met5 ;
        RECT 3458.035 1616.000 3482.985 1618.000 ;
      LAYER met5 ;
        RECT 3458.035 1599.600 3482.985 1614.400 ;
      LAYER met5 ;
        RECT 3458.035 1596.000 3482.985 1598.000 ;
      LAYER met5 ;
        RECT 3458.035 1579.600 3482.985 1594.400 ;
      LAYER met5 ;
        RECT 3458.035 1576.000 3482.985 1578.000 ;
      LAYER met5 ;
        RECT 3458.035 1559.600 3482.985 1574.400 ;
      LAYER met5 ;
        RECT 3458.035 1556.000 3482.985 1558.000 ;
      LAYER met5 ;
        RECT 3458.035 1539.600 3482.985 1554.400 ;
      LAYER met5 ;
        RECT 3458.035 1536.000 3482.985 1538.000 ;
      LAYER met5 ;
        RECT 3458.035 1519.600 3482.985 1534.400 ;
      LAYER met5 ;
        RECT 3458.035 1516.000 3482.985 1518.000 ;
      LAYER met5 ;
        RECT 3458.035 1499.600 3482.985 1514.400 ;
      LAYER met5 ;
        RECT 3458.035 1496.000 3482.985 1498.000 ;
      LAYER met5 ;
        RECT 3458.035 1479.600 3482.985 1494.400 ;
      LAYER met5 ;
        RECT 3458.035 1476.000 3482.985 1478.000 ;
      LAYER met5 ;
        RECT 3458.035 1459.600 3482.985 1474.400 ;
      LAYER met5 ;
        RECT 3458.035 1456.000 3482.985 1458.000 ;
      LAYER met5 ;
        RECT 3458.035 1439.600 3482.985 1454.400 ;
      LAYER met5 ;
        RECT 3458.035 1436.000 3482.985 1438.000 ;
      LAYER met5 ;
        RECT 3458.035 1419.600 3482.985 1434.400 ;
      LAYER met5 ;
        RECT 3458.035 1415.730 3482.985 1418.000 ;
        RECT 3563.785 1417.000 3588.000 1945.000 ;
      LAYER met5 ;
        RECT 3403.035 1414.130 3406.285 1414.435 ;
        RECT 3484.585 1414.130 3588.000 1417.000 ;
        RECT 0.000 1343.870 197.865 1350.600 ;
        RECT 3390.135 1407.400 3588.000 1414.130 ;
        RECT 0.000 1341.000 103.415 1343.870 ;
        RECT 181.715 1343.565 184.965 1343.870 ;
      LAYER met5 ;
        RECT 0.000 812.000 24.215 1341.000 ;
        RECT 105.015 1336.000 129.965 1342.270 ;
        RECT 105.015 1331.000 129.965 1333.000 ;
      LAYER met5 ;
        RECT 105.015 1314.600 129.965 1329.400 ;
      LAYER met5 ;
        RECT 105.015 1311.000 129.965 1313.000 ;
      LAYER met5 ;
        RECT 105.015 1294.600 129.965 1309.400 ;
      LAYER met5 ;
        RECT 105.015 1291.000 129.965 1293.000 ;
      LAYER met5 ;
        RECT 105.015 1274.600 129.965 1289.400 ;
      LAYER met5 ;
        RECT 105.015 1271.000 129.965 1273.000 ;
      LAYER met5 ;
        RECT 105.015 1254.600 129.965 1269.400 ;
      LAYER met5 ;
        RECT 105.015 1251.000 129.965 1253.000 ;
      LAYER met5 ;
        RECT 105.015 1234.600 129.965 1249.400 ;
      LAYER met5 ;
        RECT 105.015 1231.000 129.965 1233.000 ;
      LAYER met5 ;
        RECT 105.015 1214.600 129.965 1229.400 ;
      LAYER met5 ;
        RECT 105.015 1211.000 129.965 1213.000 ;
      LAYER met5 ;
        RECT 105.015 1194.600 129.965 1209.400 ;
      LAYER met5 ;
        RECT 105.015 1191.000 129.965 1193.000 ;
      LAYER met5 ;
        RECT 105.015 1174.600 129.965 1189.400 ;
      LAYER met5 ;
        RECT 105.015 1171.000 129.965 1173.000 ;
      LAYER met5 ;
        RECT 105.015 1154.600 129.965 1169.400 ;
      LAYER met5 ;
        RECT 105.015 1151.000 129.965 1153.000 ;
      LAYER met5 ;
        RECT 105.015 1134.600 129.965 1149.400 ;
      LAYER met5 ;
        RECT 105.015 1131.000 129.965 1133.000 ;
      LAYER met5 ;
        RECT 105.015 1114.600 129.965 1129.400 ;
      LAYER met5 ;
        RECT 105.015 1111.000 129.965 1113.000 ;
      LAYER met5 ;
        RECT 105.015 1094.600 129.965 1109.400 ;
      LAYER met5 ;
        RECT 105.015 1091.000 129.965 1093.000 ;
      LAYER met5 ;
        RECT 105.015 1074.600 129.965 1089.400 ;
      LAYER met5 ;
        RECT 105.015 1071.000 129.965 1073.000 ;
      LAYER met5 ;
        RECT 105.015 1054.600 129.965 1069.400 ;
      LAYER met5 ;
        RECT 105.015 1051.000 129.965 1053.000 ;
      LAYER met5 ;
        RECT 105.015 1034.600 129.965 1049.400 ;
      LAYER met5 ;
        RECT 105.015 1031.000 129.965 1033.000 ;
      LAYER met5 ;
        RECT 105.015 1014.600 129.965 1029.400 ;
      LAYER met5 ;
        RECT 105.015 1011.000 129.965 1013.000 ;
      LAYER met5 ;
        RECT 105.015 994.600 129.965 1009.400 ;
      LAYER met5 ;
        RECT 105.015 991.000 129.965 993.000 ;
      LAYER met5 ;
        RECT 105.015 974.600 129.965 989.400 ;
      LAYER met5 ;
        RECT 105.015 971.000 129.965 973.000 ;
      LAYER met5 ;
        RECT 105.015 954.600 129.965 969.400 ;
      LAYER met5 ;
        RECT 105.015 951.000 129.965 953.000 ;
      LAYER met5 ;
        RECT 105.015 934.600 129.965 949.400 ;
      LAYER met5 ;
        RECT 105.015 931.000 129.965 933.000 ;
      LAYER met5 ;
        RECT 105.015 914.600 129.965 929.400 ;
      LAYER met5 ;
        RECT 105.015 911.000 129.965 913.000 ;
      LAYER met5 ;
        RECT 105.015 894.600 129.965 909.400 ;
      LAYER met5 ;
        RECT 105.015 891.000 129.965 893.000 ;
      LAYER met5 ;
        RECT 105.015 874.600 129.965 889.400 ;
      LAYER met5 ;
        RECT 105.015 871.000 129.965 873.000 ;
      LAYER met5 ;
        RECT 105.015 854.600 129.965 869.400 ;
      LAYER met5 ;
        RECT 105.015 851.000 129.965 853.000 ;
      LAYER met5 ;
        RECT 105.015 834.600 129.965 849.400 ;
      LAYER met5 ;
        RECT 105.015 831.000 129.965 833.000 ;
      LAYER met5 ;
        RECT 105.015 814.600 129.965 829.400 ;
        RECT 0.000 809.130 103.415 812.000 ;
      LAYER met5 ;
        RECT 105.015 810.730 129.965 813.000 ;
        RECT 131.565 810.730 135.815 1342.270 ;
        RECT 137.415 810.730 141.665 1342.270 ;
        RECT 143.265 810.730 152.265 1342.270 ;
        RECT 153.865 810.730 158.315 1342.270 ;
        RECT 159.915 1341.000 163.160 1342.270 ;
        RECT 159.915 812.000 163.165 1341.000 ;
        RECT 159.915 810.730 163.160 812.000 ;
        RECT 164.765 810.730 168.015 1342.270 ;
        RECT 169.615 810.730 174.065 1342.270 ;
        RECT 175.665 810.730 180.115 1342.270 ;
        RECT 181.715 810.970 184.965 1341.965 ;
        RECT 186.565 810.730 191.015 1342.270 ;
        RECT 192.615 810.730 197.865 1342.270 ;
      LAYER met5 ;
        RECT 3390.135 1341.600 3490.960 1407.400 ;
        RECT 3556.610 1341.600 3588.000 1407.400 ;
        RECT 3390.135 1339.870 3588.000 1341.600 ;
        RECT 3403.035 1339.630 3406.285 1339.870 ;
        RECT 181.715 809.130 184.965 809.370 ;
        RECT 0.000 807.400 197.865 809.130 ;
        RECT 0.000 741.600 31.390 807.400 ;
        RECT 97.040 741.600 197.865 807.400 ;
      LAYER met5 ;
        RECT 3390.135 806.730 3395.385 1338.270 ;
        RECT 3396.985 806.730 3401.435 1338.270 ;
        RECT 3403.035 807.035 3406.285 1338.030 ;
        RECT 3407.885 806.730 3412.335 1338.270 ;
        RECT 3413.935 806.730 3418.385 1338.270 ;
        RECT 3419.985 806.730 3423.235 1338.270 ;
        RECT 3424.840 1337.000 3428.085 1338.270 ;
        RECT 3424.835 808.000 3428.085 1337.000 ;
        RECT 3424.840 806.730 3428.085 808.000 ;
        RECT 3429.685 806.730 3434.135 1338.270 ;
        RECT 3435.735 806.730 3444.735 1338.270 ;
        RECT 3446.335 806.730 3450.585 1338.270 ;
        RECT 3452.185 806.730 3456.435 1338.270 ;
        RECT 3458.035 1332.000 3482.985 1338.270 ;
      LAYER met5 ;
        RECT 3484.585 1337.000 3588.000 1339.870 ;
      LAYER met5 ;
        RECT 3458.035 1327.000 3482.985 1329.000 ;
      LAYER met5 ;
        RECT 3458.035 1310.600 3482.985 1325.400 ;
      LAYER met5 ;
        RECT 3458.035 1307.000 3482.985 1309.000 ;
      LAYER met5 ;
        RECT 3458.035 1290.600 3482.985 1305.400 ;
      LAYER met5 ;
        RECT 3458.035 1287.000 3482.985 1289.000 ;
      LAYER met5 ;
        RECT 3458.035 1270.600 3482.985 1285.400 ;
      LAYER met5 ;
        RECT 3458.035 1267.000 3482.985 1269.000 ;
      LAYER met5 ;
        RECT 3458.035 1250.600 3482.985 1265.400 ;
      LAYER met5 ;
        RECT 3458.035 1247.000 3482.985 1249.000 ;
      LAYER met5 ;
        RECT 3458.035 1230.600 3482.985 1245.400 ;
      LAYER met5 ;
        RECT 3458.035 1227.000 3482.985 1229.000 ;
      LAYER met5 ;
        RECT 3458.035 1210.600 3482.985 1225.400 ;
      LAYER met5 ;
        RECT 3458.035 1207.000 3482.985 1209.000 ;
      LAYER met5 ;
        RECT 3458.035 1190.600 3482.985 1205.400 ;
      LAYER met5 ;
        RECT 3458.035 1187.000 3482.985 1189.000 ;
      LAYER met5 ;
        RECT 3458.035 1170.600 3482.985 1185.400 ;
      LAYER met5 ;
        RECT 3458.035 1167.000 3482.985 1169.000 ;
      LAYER met5 ;
        RECT 3458.035 1150.600 3482.985 1165.400 ;
      LAYER met5 ;
        RECT 3458.035 1147.000 3482.985 1149.000 ;
      LAYER met5 ;
        RECT 3458.035 1130.600 3482.985 1145.400 ;
      LAYER met5 ;
        RECT 3458.035 1127.000 3482.985 1129.000 ;
      LAYER met5 ;
        RECT 3458.035 1110.600 3482.985 1125.400 ;
      LAYER met5 ;
        RECT 3458.035 1107.000 3482.985 1109.000 ;
      LAYER met5 ;
        RECT 3458.035 1090.600 3482.985 1105.400 ;
      LAYER met5 ;
        RECT 3458.035 1087.000 3482.985 1089.000 ;
      LAYER met5 ;
        RECT 3458.035 1070.600 3482.985 1085.400 ;
      LAYER met5 ;
        RECT 3458.035 1067.000 3482.985 1069.000 ;
      LAYER met5 ;
        RECT 3458.035 1050.600 3482.985 1065.400 ;
      LAYER met5 ;
        RECT 3458.035 1047.000 3482.985 1049.000 ;
      LAYER met5 ;
        RECT 3458.035 1030.600 3482.985 1045.400 ;
      LAYER met5 ;
        RECT 3458.035 1027.000 3482.985 1029.000 ;
      LAYER met5 ;
        RECT 3458.035 1010.600 3482.985 1025.400 ;
      LAYER met5 ;
        RECT 3458.035 1007.000 3482.985 1009.000 ;
      LAYER met5 ;
        RECT 3458.035 990.600 3482.985 1005.400 ;
      LAYER met5 ;
        RECT 3458.035 987.000 3482.985 989.000 ;
      LAYER met5 ;
        RECT 3458.035 970.600 3482.985 985.400 ;
      LAYER met5 ;
        RECT 3458.035 967.000 3482.985 969.000 ;
      LAYER met5 ;
        RECT 3458.035 950.600 3482.985 965.400 ;
      LAYER met5 ;
        RECT 3458.035 947.000 3482.985 949.000 ;
      LAYER met5 ;
        RECT 3458.035 930.600 3482.985 945.400 ;
      LAYER met5 ;
        RECT 3458.035 927.000 3482.985 929.000 ;
      LAYER met5 ;
        RECT 3458.035 910.600 3482.985 925.400 ;
      LAYER met5 ;
        RECT 3458.035 907.000 3482.985 909.000 ;
      LAYER met5 ;
        RECT 3458.035 890.600 3482.985 905.400 ;
      LAYER met5 ;
        RECT 3458.035 887.000 3482.985 889.000 ;
      LAYER met5 ;
        RECT 3458.035 870.600 3482.985 885.400 ;
      LAYER met5 ;
        RECT 3458.035 867.000 3482.985 869.000 ;
      LAYER met5 ;
        RECT 3458.035 850.600 3482.985 865.400 ;
      LAYER met5 ;
        RECT 3458.035 847.000 3482.985 849.000 ;
      LAYER met5 ;
        RECT 3458.035 830.600 3482.985 845.400 ;
      LAYER met5 ;
        RECT 3458.035 827.000 3482.985 829.000 ;
      LAYER met5 ;
        RECT 3458.035 810.600 3482.985 825.400 ;
      LAYER met5 ;
        RECT 3458.035 806.730 3482.985 809.000 ;
        RECT 3563.785 808.000 3588.000 1337.000 ;
      LAYER met5 ;
        RECT 3403.035 805.130 3406.285 805.435 ;
        RECT 3484.585 805.130 3588.000 808.000 ;
        RECT 0.000 734.870 197.865 741.600 ;
        RECT 3390.135 798.400 3588.000 805.130 ;
        RECT 0.000 732.000 103.415 734.870 ;
        RECT 181.715 734.565 184.965 734.870 ;
      LAYER met5 ;
        RECT 0.000 204.000 24.215 732.000 ;
        RECT 105.015 728.000 129.965 733.270 ;
        RECT 105.015 723.000 129.965 725.000 ;
      LAYER met5 ;
        RECT 105.015 706.600 129.965 721.400 ;
      LAYER met5 ;
        RECT 105.015 703.000 129.965 705.000 ;
      LAYER met5 ;
        RECT 105.015 686.600 129.965 701.400 ;
      LAYER met5 ;
        RECT 105.015 683.000 129.965 685.000 ;
      LAYER met5 ;
        RECT 105.015 666.600 129.965 681.400 ;
      LAYER met5 ;
        RECT 105.015 663.000 129.965 665.000 ;
      LAYER met5 ;
        RECT 105.015 646.600 129.965 661.400 ;
      LAYER met5 ;
        RECT 105.015 643.000 129.965 645.000 ;
      LAYER met5 ;
        RECT 105.015 626.600 129.965 641.400 ;
      LAYER met5 ;
        RECT 105.015 623.000 129.965 625.000 ;
      LAYER met5 ;
        RECT 105.015 606.600 129.965 621.400 ;
      LAYER met5 ;
        RECT 105.015 603.000 129.965 605.000 ;
      LAYER met5 ;
        RECT 105.015 586.600 129.965 601.400 ;
      LAYER met5 ;
        RECT 105.015 583.000 129.965 585.000 ;
      LAYER met5 ;
        RECT 105.015 566.600 129.965 581.400 ;
      LAYER met5 ;
        RECT 105.015 563.000 129.965 565.000 ;
      LAYER met5 ;
        RECT 105.015 546.600 129.965 561.400 ;
      LAYER met5 ;
        RECT 105.015 543.000 129.965 545.000 ;
      LAYER met5 ;
        RECT 105.015 526.600 129.965 541.400 ;
      LAYER met5 ;
        RECT 105.015 523.000 129.965 525.000 ;
      LAYER met5 ;
        RECT 105.015 506.600 129.965 521.400 ;
      LAYER met5 ;
        RECT 105.015 503.000 129.965 505.000 ;
      LAYER met5 ;
        RECT 105.015 486.600 129.965 501.400 ;
      LAYER met5 ;
        RECT 105.015 483.000 129.965 485.000 ;
      LAYER met5 ;
        RECT 105.015 466.600 129.965 481.400 ;
      LAYER met5 ;
        RECT 105.015 463.000 129.965 465.000 ;
      LAYER met5 ;
        RECT 105.015 446.600 129.965 461.400 ;
      LAYER met5 ;
        RECT 105.015 443.000 129.965 445.000 ;
      LAYER met5 ;
        RECT 105.015 426.600 129.965 441.400 ;
      LAYER met5 ;
        RECT 105.015 423.000 129.965 425.000 ;
      LAYER met5 ;
        RECT 105.015 406.600 129.965 421.400 ;
      LAYER met5 ;
        RECT 105.015 403.000 129.965 405.000 ;
      LAYER met5 ;
        RECT 105.015 386.600 129.965 401.400 ;
      LAYER met5 ;
        RECT 105.015 383.000 129.965 385.000 ;
      LAYER met5 ;
        RECT 105.015 366.600 129.965 381.400 ;
      LAYER met5 ;
        RECT 105.015 363.000 129.965 365.000 ;
      LAYER met5 ;
        RECT 105.015 346.600 129.965 361.400 ;
      LAYER met5 ;
        RECT 105.015 343.000 129.965 345.000 ;
      LAYER met5 ;
        RECT 105.015 326.600 129.965 341.400 ;
      LAYER met5 ;
        RECT 105.015 323.000 129.965 325.000 ;
      LAYER met5 ;
        RECT 105.015 306.600 129.965 321.400 ;
      LAYER met5 ;
        RECT 105.015 303.000 129.965 305.000 ;
      LAYER met5 ;
        RECT 105.015 286.600 129.965 301.400 ;
      LAYER met5 ;
        RECT 105.015 283.000 129.965 285.000 ;
      LAYER met5 ;
        RECT 105.015 266.600 129.965 281.400 ;
      LAYER met5 ;
        RECT 105.015 263.000 129.965 265.000 ;
      LAYER met5 ;
        RECT 105.015 246.600 129.965 261.400 ;
      LAYER met5 ;
        RECT 105.015 243.000 129.965 245.000 ;
      LAYER met5 ;
        RECT 105.015 226.600 129.965 241.400 ;
      LAYER met5 ;
        RECT 105.015 223.000 129.965 225.000 ;
      LAYER met5 ;
        RECT 105.015 206.600 129.965 221.400 ;
        RECT 0.000 200.545 103.415 204.000 ;
      LAYER met5 ;
        RECT 105.015 202.145 129.965 205.000 ;
        RECT 131.565 202.730 135.815 733.270 ;
        RECT 137.415 202.730 141.665 733.270 ;
      LAYER met5 ;
        RECT 131.565 200.545 141.665 201.130 ;
        RECT 0.000 175.245 141.665 200.545 ;
      LAYER met5 ;
        RECT 143.265 176.845 152.265 733.270 ;
        RECT 153.865 202.730 158.315 733.270 ;
        RECT 159.915 732.000 163.160 733.270 ;
        RECT 159.915 204.000 163.165 732.000 ;
        RECT 159.915 202.730 163.160 204.000 ;
        RECT 164.765 202.730 168.015 733.270 ;
        RECT 169.615 202.730 174.065 733.270 ;
        RECT 175.665 202.730 180.115 733.270 ;
        RECT 181.715 202.745 184.965 732.965 ;
        RECT 186.565 202.730 191.015 733.270 ;
        RECT 192.615 202.730 197.865 733.270 ;
      LAYER met5 ;
        RECT 3390.135 732.600 3490.960 798.400 ;
        RECT 3556.610 732.600 3588.000 798.400 ;
        RECT 3390.135 730.870 3588.000 732.600 ;
        RECT 3403.035 730.630 3406.285 730.870 ;
        RECT 181.715 201.130 184.965 201.145 ;
        RECT 199.465 201.130 200.000 204.000 ;
        RECT 153.865 199.465 200.000 201.130 ;
        RECT 3384.000 199.465 3388.535 200.000 ;
        RECT 153.865 192.615 196.050 199.465 ;
      LAYER met5 ;
        RECT 197.650 192.615 668.270 197.865 ;
      LAYER met5 ;
        RECT 153.865 184.965 194.615 192.615 ;
      LAYER met5 ;
        RECT 196.215 186.565 668.270 191.015 ;
      LAYER met5 ;
        RECT 669.870 184.965 739.130 197.865 ;
      LAYER met5 ;
        RECT 740.730 192.615 1210.270 197.865 ;
        RECT 740.730 186.565 1210.270 191.015 ;
      LAYER met5 ;
        RECT 1211.870 184.965 1284.000 197.865 ;
      LAYER met5 ;
        RECT 1284.000 192.615 1753.270 197.865 ;
        RECT 1284.000 186.565 1753.270 191.015 ;
      LAYER met5 ;
        RECT 1754.870 184.965 1829.130 197.865 ;
      LAYER met5 ;
        RECT 1830.730 192.615 2300.270 197.865 ;
        RECT 1830.730 186.565 2300.270 191.015 ;
      LAYER met5 ;
        RECT 2301.870 184.965 2371.130 197.865 ;
      LAYER met5 ;
        RECT 2372.730 192.615 2842.270 197.865 ;
        RECT 2372.730 186.565 2842.270 191.015 ;
      LAYER met5 ;
        RECT 2843.870 184.965 2913.130 197.865 ;
      LAYER met5 ;
        RECT 2914.730 192.615 3385.270 197.865 ;
      LAYER met5 ;
        RECT 3386.870 196.050 3388.535 199.465 ;
      LAYER met5 ;
        RECT 3390.135 197.650 3395.385 729.270 ;
        RECT 3396.985 196.215 3401.435 729.270 ;
        RECT 3403.035 198.530 3406.285 729.030 ;
        RECT 3407.885 198.475 3412.335 729.270 ;
        RECT 3413.935 198.400 3418.385 729.270 ;
        RECT 3419.985 198.615 3423.235 729.270 ;
        RECT 3424.840 728.000 3428.085 729.270 ;
        RECT 3424.835 198.665 3428.085 728.000 ;
        RECT 3429.685 198.525 3434.135 729.270 ;
      LAYER met5 ;
        RECT 3424.835 197.015 3428.085 197.065 ;
        RECT 3403.035 196.875 3406.285 196.930 ;
        RECT 3419.985 196.925 3428.085 197.015 ;
        RECT 3403.035 196.800 3412.335 196.875 ;
        RECT 3419.985 196.800 3434.135 196.925 ;
        RECT 3386.870 194.615 3395.385 196.050 ;
        RECT 3403.035 194.615 3434.135 196.800 ;
      LAYER met5 ;
        RECT 2914.730 186.565 3385.270 191.015 ;
      LAYER met5 ;
        RECT 3386.870 184.965 3434.135 194.615 ;
        RECT 153.865 181.715 196.930 184.965 ;
      LAYER met5 ;
        RECT 198.530 181.715 667.965 184.965 ;
      LAYER met5 ;
        RECT 669.565 181.715 739.435 184.965 ;
      LAYER met5 ;
        RECT 741.035 181.715 1209.965 184.965 ;
      LAYER met5 ;
        RECT 153.865 175.665 196.875 181.715 ;
      LAYER met5 ;
        RECT 198.475 175.665 668.270 180.115 ;
      LAYER met5 ;
        RECT 153.865 175.245 196.800 175.665 ;
        RECT 0.000 168.015 196.800 175.245 ;
      LAYER met5 ;
        RECT 198.400 169.615 668.270 174.065 ;
      LAYER met5 ;
        RECT 0.000 163.165 197.015 168.015 ;
      LAYER met5 ;
        RECT 198.615 164.765 668.270 168.015 ;
      LAYER met5 ;
        RECT 0.000 159.915 197.065 163.165 ;
      LAYER met5 ;
        RECT 198.665 163.160 667.000 163.165 ;
        RECT 198.665 159.915 668.270 163.160 ;
      LAYER met5 ;
        RECT 0.000 153.865 196.925 159.915 ;
      LAYER met5 ;
        RECT 198.525 153.865 668.270 158.315 ;
      LAYER met5 ;
        RECT 0.000 141.665 175.245 153.865 ;
      LAYER met5 ;
        RECT 176.845 143.265 668.270 152.265 ;
      LAYER met5 ;
        RECT 0.000 135.815 196.775 141.665 ;
      LAYER met5 ;
        RECT 198.375 137.415 668.270 141.665 ;
      LAYER met5 ;
        RECT 0.000 131.565 196.920 135.815 ;
      LAYER met5 ;
        RECT 198.520 131.565 668.270 135.815 ;
      LAYER met5 ;
        RECT 0.000 103.415 195.755 131.565 ;
      LAYER met5 ;
        RECT 197.355 105.015 201.000 129.965 ;
      LAYER met5 ;
        RECT 202.600 105.015 217.400 129.965 ;
      LAYER met5 ;
        RECT 219.000 105.015 221.000 129.965 ;
      LAYER met5 ;
        RECT 222.600 105.015 237.400 129.965 ;
      LAYER met5 ;
        RECT 239.000 105.015 241.000 129.965 ;
      LAYER met5 ;
        RECT 242.600 105.015 257.400 129.965 ;
      LAYER met5 ;
        RECT 259.000 105.015 261.000 129.965 ;
      LAYER met5 ;
        RECT 262.600 105.015 277.400 129.965 ;
      LAYER met5 ;
        RECT 279.000 105.015 281.000 129.965 ;
      LAYER met5 ;
        RECT 282.600 105.015 297.400 129.965 ;
      LAYER met5 ;
        RECT 299.000 105.015 301.000 129.965 ;
      LAYER met5 ;
        RECT 302.600 105.015 317.400 129.965 ;
      LAYER met5 ;
        RECT 319.000 105.015 321.000 129.965 ;
      LAYER met5 ;
        RECT 322.600 105.015 337.400 129.965 ;
      LAYER met5 ;
        RECT 339.000 105.015 341.000 129.965 ;
      LAYER met5 ;
        RECT 342.600 105.015 357.400 129.965 ;
      LAYER met5 ;
        RECT 359.000 105.015 361.000 129.965 ;
      LAYER met5 ;
        RECT 362.600 105.015 377.400 129.965 ;
      LAYER met5 ;
        RECT 379.000 105.015 381.000 129.965 ;
      LAYER met5 ;
        RECT 382.600 105.015 397.400 129.965 ;
      LAYER met5 ;
        RECT 399.000 105.015 401.000 129.965 ;
      LAYER met5 ;
        RECT 402.600 105.015 417.400 129.965 ;
      LAYER met5 ;
        RECT 419.000 105.015 421.000 129.965 ;
      LAYER met5 ;
        RECT 422.600 105.015 437.400 129.965 ;
      LAYER met5 ;
        RECT 439.000 105.015 441.000 129.965 ;
      LAYER met5 ;
        RECT 442.600 105.015 457.400 129.965 ;
      LAYER met5 ;
        RECT 459.000 105.015 461.000 129.965 ;
      LAYER met5 ;
        RECT 462.600 105.015 477.400 129.965 ;
      LAYER met5 ;
        RECT 479.000 105.015 481.000 129.965 ;
      LAYER met5 ;
        RECT 482.600 105.015 497.400 129.965 ;
      LAYER met5 ;
        RECT 499.000 105.015 501.000 129.965 ;
      LAYER met5 ;
        RECT 502.600 105.015 517.400 129.965 ;
      LAYER met5 ;
        RECT 519.000 105.015 521.000 129.965 ;
      LAYER met5 ;
        RECT 522.600 105.015 537.400 129.965 ;
      LAYER met5 ;
        RECT 539.000 105.015 541.000 129.965 ;
      LAYER met5 ;
        RECT 542.600 105.015 557.400 129.965 ;
      LAYER met5 ;
        RECT 559.000 105.015 561.000 129.965 ;
      LAYER met5 ;
        RECT 562.600 105.015 577.400 129.965 ;
      LAYER met5 ;
        RECT 579.000 105.015 581.000 129.965 ;
      LAYER met5 ;
        RECT 582.600 105.015 597.400 129.965 ;
      LAYER met5 ;
        RECT 599.000 105.015 601.000 129.965 ;
      LAYER met5 ;
        RECT 602.600 105.015 617.400 129.965 ;
      LAYER met5 ;
        RECT 619.000 105.015 621.000 129.965 ;
      LAYER met5 ;
        RECT 622.600 105.015 637.400 129.965 ;
      LAYER met5 ;
        RECT 639.000 105.015 641.000 129.965 ;
      LAYER met5 ;
        RECT 642.600 105.015 657.400 129.965 ;
      LAYER met5 ;
        RECT 659.000 105.015 661.000 129.965 ;
        RECT 664.000 105.015 668.270 129.965 ;
      LAYER met5 ;
        RECT 669.870 103.415 739.130 181.715 ;
        RECT 1211.565 180.115 1284.000 184.965 ;
      LAYER met5 ;
        RECT 1284.000 181.715 1753.030 184.965 ;
      LAYER met5 ;
        RECT 1754.630 181.715 1829.435 184.965 ;
      LAYER met5 ;
        RECT 1831.035 181.715 2299.965 184.965 ;
      LAYER met5 ;
        RECT 2301.565 181.715 2371.435 184.965 ;
      LAYER met5 ;
        RECT 2373.035 181.715 2841.965 184.965 ;
      LAYER met5 ;
        RECT 2843.565 181.715 2913.435 184.965 ;
      LAYER met5 ;
        RECT 2915.035 181.715 3385.255 184.965 ;
      LAYER met5 ;
        RECT 3386.855 181.715 3434.135 184.965 ;
      LAYER met5 ;
        RECT 740.730 175.665 1209.000 180.115 ;
      LAYER met5 ;
        RECT 1209.000 175.665 1284.000 180.115 ;
      LAYER met5 ;
        RECT 1284.000 175.665 1753.270 180.115 ;
        RECT 740.730 169.615 1210.270 174.065 ;
        RECT 740.730 164.765 1210.270 168.015 ;
      LAYER met5 ;
        RECT 1211.870 163.165 1284.000 175.665 ;
      LAYER met5 ;
        RECT 1284.000 169.615 1753.270 174.065 ;
        RECT 1284.000 164.765 1753.270 168.015 ;
        RECT 742.000 163.160 1209.000 163.165 ;
        RECT 740.730 159.915 1209.000 163.160 ;
      LAYER met5 ;
        RECT 1209.000 159.915 1284.000 163.165 ;
      LAYER met5 ;
        RECT 1284.000 163.160 1752.000 163.165 ;
        RECT 1284.000 159.915 1753.270 163.160 ;
        RECT 740.730 153.865 1210.270 158.315 ;
        RECT 740.730 143.265 1210.270 152.265 ;
        RECT 740.730 137.415 1210.270 141.665 ;
        RECT 740.730 131.565 1210.270 135.815 ;
        RECT 740.730 105.015 743.000 129.965 ;
      LAYER met5 ;
        RECT 744.600 105.015 759.400 129.965 ;
      LAYER met5 ;
        RECT 761.000 105.015 763.000 129.965 ;
      LAYER met5 ;
        RECT 764.600 105.015 779.400 129.965 ;
      LAYER met5 ;
        RECT 781.000 105.015 783.000 129.965 ;
      LAYER met5 ;
        RECT 784.600 105.015 799.400 129.965 ;
      LAYER met5 ;
        RECT 801.000 105.015 803.000 129.965 ;
      LAYER met5 ;
        RECT 804.600 105.015 819.400 129.965 ;
      LAYER met5 ;
        RECT 821.000 105.015 823.000 129.965 ;
      LAYER met5 ;
        RECT 824.600 105.015 839.400 129.965 ;
      LAYER met5 ;
        RECT 841.000 105.015 843.000 129.965 ;
      LAYER met5 ;
        RECT 844.600 105.015 859.400 129.965 ;
      LAYER met5 ;
        RECT 861.000 105.015 863.000 129.965 ;
      LAYER met5 ;
        RECT 864.600 105.015 879.400 129.965 ;
      LAYER met5 ;
        RECT 881.000 105.015 883.000 129.965 ;
      LAYER met5 ;
        RECT 884.600 105.015 899.400 129.965 ;
      LAYER met5 ;
        RECT 901.000 105.015 903.000 129.965 ;
      LAYER met5 ;
        RECT 904.600 105.015 919.400 129.965 ;
      LAYER met5 ;
        RECT 921.000 105.015 923.000 129.965 ;
      LAYER met5 ;
        RECT 924.600 105.015 939.400 129.965 ;
      LAYER met5 ;
        RECT 941.000 105.015 943.000 129.965 ;
      LAYER met5 ;
        RECT 944.600 105.015 959.400 129.965 ;
      LAYER met5 ;
        RECT 961.000 105.015 963.000 129.965 ;
      LAYER met5 ;
        RECT 964.600 105.015 979.400 129.965 ;
      LAYER met5 ;
        RECT 981.000 105.015 983.000 129.965 ;
      LAYER met5 ;
        RECT 984.600 105.015 999.400 129.965 ;
      LAYER met5 ;
        RECT 1001.000 105.015 1003.000 129.965 ;
      LAYER met5 ;
        RECT 1004.600 105.015 1019.400 129.965 ;
      LAYER met5 ;
        RECT 1021.000 105.015 1023.000 129.965 ;
      LAYER met5 ;
        RECT 1024.600 105.015 1039.400 129.965 ;
      LAYER met5 ;
        RECT 1041.000 105.015 1043.000 129.965 ;
      LAYER met5 ;
        RECT 1044.600 105.015 1059.400 129.965 ;
      LAYER met5 ;
        RECT 1061.000 105.015 1063.000 129.965 ;
      LAYER met5 ;
        RECT 1064.600 105.015 1079.400 129.965 ;
      LAYER met5 ;
        RECT 1081.000 105.015 1083.000 129.965 ;
      LAYER met5 ;
        RECT 1084.600 105.015 1099.400 129.965 ;
      LAYER met5 ;
        RECT 1101.000 105.015 1103.000 129.965 ;
      LAYER met5 ;
        RECT 1104.600 105.015 1119.400 129.965 ;
      LAYER met5 ;
        RECT 1121.000 105.015 1123.000 129.965 ;
      LAYER met5 ;
        RECT 1124.600 105.015 1139.400 129.965 ;
      LAYER met5 ;
        RECT 1141.000 105.015 1143.000 129.965 ;
      LAYER met5 ;
        RECT 1144.600 105.015 1159.400 129.965 ;
      LAYER met5 ;
        RECT 1161.000 105.015 1163.000 129.965 ;
      LAYER met5 ;
        RECT 1164.600 105.015 1179.400 129.965 ;
      LAYER met5 ;
        RECT 1181.000 105.015 1183.000 129.965 ;
      LAYER met5 ;
        RECT 1184.600 105.015 1199.400 129.965 ;
      LAYER met5 ;
        RECT 1201.000 105.015 1203.000 129.965 ;
        RECT 1206.000 105.015 1210.270 129.965 ;
      LAYER met5 ;
        RECT 1211.870 103.415 1284.000 159.915 ;
      LAYER met5 ;
        RECT 1284.000 153.865 1753.270 158.315 ;
        RECT 1284.000 143.265 1753.270 152.265 ;
        RECT 1284.000 137.415 1753.270 141.665 ;
        RECT 1284.000 131.565 1753.270 135.815 ;
        RECT 1284.000 105.015 1285.000 129.965 ;
      LAYER met5 ;
        RECT 1286.600 105.015 1301.400 129.965 ;
      LAYER met5 ;
        RECT 1303.000 105.015 1305.000 129.965 ;
      LAYER met5 ;
        RECT 1306.600 105.015 1321.400 129.965 ;
      LAYER met5 ;
        RECT 1323.000 105.015 1325.000 129.965 ;
      LAYER met5 ;
        RECT 1326.600 105.015 1341.400 129.965 ;
      LAYER met5 ;
        RECT 1343.000 105.015 1345.000 129.965 ;
      LAYER met5 ;
        RECT 1346.600 105.015 1361.400 129.965 ;
      LAYER met5 ;
        RECT 1363.000 105.015 1365.000 129.965 ;
      LAYER met5 ;
        RECT 1366.600 105.015 1381.400 129.965 ;
      LAYER met5 ;
        RECT 1383.000 105.015 1385.000 129.965 ;
      LAYER met5 ;
        RECT 1386.600 105.015 1401.400 129.965 ;
      LAYER met5 ;
        RECT 1403.000 105.015 1405.000 129.965 ;
      LAYER met5 ;
        RECT 1406.600 105.015 1421.400 129.965 ;
      LAYER met5 ;
        RECT 1423.000 105.015 1425.000 129.965 ;
      LAYER met5 ;
        RECT 1426.600 105.015 1441.400 129.965 ;
      LAYER met5 ;
        RECT 1443.000 105.015 1445.000 129.965 ;
      LAYER met5 ;
        RECT 1446.600 105.015 1461.400 129.965 ;
      LAYER met5 ;
        RECT 1463.000 105.015 1465.000 129.965 ;
      LAYER met5 ;
        RECT 1466.600 105.015 1481.400 129.965 ;
      LAYER met5 ;
        RECT 1483.000 105.015 1485.000 129.965 ;
      LAYER met5 ;
        RECT 1486.600 105.015 1501.400 129.965 ;
      LAYER met5 ;
        RECT 1503.000 105.015 1505.000 129.965 ;
      LAYER met5 ;
        RECT 1506.600 105.015 1521.400 129.965 ;
      LAYER met5 ;
        RECT 1523.000 105.015 1525.000 129.965 ;
      LAYER met5 ;
        RECT 1526.600 105.015 1541.400 129.965 ;
      LAYER met5 ;
        RECT 1543.000 105.015 1545.000 129.965 ;
      LAYER met5 ;
        RECT 1546.600 105.015 1561.400 129.965 ;
      LAYER met5 ;
        RECT 1563.000 105.015 1565.000 129.965 ;
      LAYER met5 ;
        RECT 1566.600 105.015 1581.400 129.965 ;
      LAYER met5 ;
        RECT 1583.000 105.015 1585.000 129.965 ;
      LAYER met5 ;
        RECT 1586.600 105.015 1601.400 129.965 ;
      LAYER met5 ;
        RECT 1603.000 105.015 1605.000 129.965 ;
      LAYER met5 ;
        RECT 1606.600 105.015 1621.400 129.965 ;
      LAYER met5 ;
        RECT 1623.000 105.015 1625.000 129.965 ;
      LAYER met5 ;
        RECT 1626.600 105.015 1641.400 129.965 ;
      LAYER met5 ;
        RECT 1643.000 105.015 1645.000 129.965 ;
      LAYER met5 ;
        RECT 1646.600 105.015 1661.400 129.965 ;
      LAYER met5 ;
        RECT 1663.000 105.015 1665.000 129.965 ;
      LAYER met5 ;
        RECT 1666.600 105.015 1681.400 129.965 ;
      LAYER met5 ;
        RECT 1683.000 105.015 1685.000 129.965 ;
      LAYER met5 ;
        RECT 1686.600 105.015 1701.400 129.965 ;
      LAYER met5 ;
        RECT 1703.000 105.015 1705.000 129.965 ;
      LAYER met5 ;
        RECT 1706.600 105.015 1721.400 129.965 ;
      LAYER met5 ;
        RECT 1723.000 105.015 1725.000 129.965 ;
      LAYER met5 ;
        RECT 1726.600 105.015 1741.400 129.965 ;
      LAYER met5 ;
        RECT 1743.000 105.015 1745.000 129.965 ;
        RECT 1748.000 105.015 1753.270 129.965 ;
      LAYER met5 ;
        RECT 1754.870 103.415 1829.130 181.715 ;
      LAYER met5 ;
        RECT 1830.730 175.665 2300.270 180.115 ;
        RECT 1830.730 169.615 2300.270 174.065 ;
        RECT 1830.730 164.765 2300.270 168.015 ;
        RECT 1832.000 163.160 2299.000 163.165 ;
        RECT 1830.730 159.915 2300.270 163.160 ;
        RECT 1830.730 153.865 2300.270 158.315 ;
        RECT 1830.730 143.265 2300.270 152.265 ;
        RECT 1830.730 137.415 2300.270 141.665 ;
        RECT 1830.730 131.565 2300.270 135.815 ;
        RECT 1830.730 105.015 1833.000 129.965 ;
      LAYER met5 ;
        RECT 1834.600 105.015 1849.400 129.965 ;
      LAYER met5 ;
        RECT 1851.000 105.015 1853.000 129.965 ;
      LAYER met5 ;
        RECT 1854.600 105.015 1869.400 129.965 ;
      LAYER met5 ;
        RECT 1871.000 105.015 1873.000 129.965 ;
      LAYER met5 ;
        RECT 1874.600 105.015 1889.400 129.965 ;
      LAYER met5 ;
        RECT 1891.000 105.015 1893.000 129.965 ;
      LAYER met5 ;
        RECT 1894.600 105.015 1909.400 129.965 ;
      LAYER met5 ;
        RECT 1911.000 105.015 1913.000 129.965 ;
      LAYER met5 ;
        RECT 1914.600 105.015 1929.400 129.965 ;
      LAYER met5 ;
        RECT 1931.000 105.015 1933.000 129.965 ;
      LAYER met5 ;
        RECT 1934.600 105.015 1949.400 129.965 ;
      LAYER met5 ;
        RECT 1951.000 105.015 1953.000 129.965 ;
      LAYER met5 ;
        RECT 1954.600 105.015 1969.400 129.965 ;
      LAYER met5 ;
        RECT 1971.000 105.015 1973.000 129.965 ;
      LAYER met5 ;
        RECT 1974.600 105.015 1989.400 129.965 ;
      LAYER met5 ;
        RECT 1991.000 105.015 1993.000 129.965 ;
      LAYER met5 ;
        RECT 1994.600 105.015 2009.400 129.965 ;
      LAYER met5 ;
        RECT 2011.000 105.015 2013.000 129.965 ;
      LAYER met5 ;
        RECT 2014.600 105.015 2029.400 129.965 ;
      LAYER met5 ;
        RECT 2031.000 105.015 2033.000 129.965 ;
      LAYER met5 ;
        RECT 2034.600 105.015 2049.400 129.965 ;
      LAYER met5 ;
        RECT 2051.000 105.015 2053.000 129.965 ;
      LAYER met5 ;
        RECT 2054.600 105.015 2069.400 129.965 ;
      LAYER met5 ;
        RECT 2071.000 105.015 2073.000 129.965 ;
      LAYER met5 ;
        RECT 2074.600 105.015 2089.400 129.965 ;
      LAYER met5 ;
        RECT 2091.000 105.015 2093.000 129.965 ;
      LAYER met5 ;
        RECT 2094.600 105.015 2109.400 129.965 ;
      LAYER met5 ;
        RECT 2111.000 105.015 2113.000 129.965 ;
      LAYER met5 ;
        RECT 2114.600 105.015 2129.400 129.965 ;
      LAYER met5 ;
        RECT 2131.000 105.015 2133.000 129.965 ;
      LAYER met5 ;
        RECT 2134.600 105.015 2149.400 129.965 ;
      LAYER met5 ;
        RECT 2151.000 105.015 2153.000 129.965 ;
      LAYER met5 ;
        RECT 2154.600 105.015 2169.400 129.965 ;
      LAYER met5 ;
        RECT 2171.000 105.015 2173.000 129.965 ;
      LAYER met5 ;
        RECT 2174.600 105.015 2189.400 129.965 ;
      LAYER met5 ;
        RECT 2191.000 105.015 2193.000 129.965 ;
      LAYER met5 ;
        RECT 2194.600 105.015 2209.400 129.965 ;
      LAYER met5 ;
        RECT 2211.000 105.015 2213.000 129.965 ;
      LAYER met5 ;
        RECT 2214.600 105.015 2229.400 129.965 ;
      LAYER met5 ;
        RECT 2231.000 105.015 2233.000 129.965 ;
      LAYER met5 ;
        RECT 2234.600 105.015 2249.400 129.965 ;
      LAYER met5 ;
        RECT 2251.000 105.015 2253.000 129.965 ;
      LAYER met5 ;
        RECT 2254.600 105.015 2269.400 129.965 ;
      LAYER met5 ;
        RECT 2271.000 105.015 2273.000 129.965 ;
      LAYER met5 ;
        RECT 2274.600 105.015 2289.400 129.965 ;
      LAYER met5 ;
        RECT 2291.000 105.015 2293.000 129.965 ;
        RECT 2296.000 105.015 2300.270 129.965 ;
      LAYER met5 ;
        RECT 2301.870 103.415 2371.130 181.715 ;
      LAYER met5 ;
        RECT 2372.730 175.665 2842.270 180.115 ;
        RECT 2372.730 169.615 2842.270 174.065 ;
        RECT 2372.730 164.765 2842.270 168.015 ;
        RECT 2374.000 163.160 2841.000 163.165 ;
        RECT 2372.730 159.915 2842.270 163.160 ;
        RECT 2372.730 153.865 2842.270 158.315 ;
        RECT 2372.730 143.265 2842.270 152.265 ;
        RECT 2372.730 137.415 2842.270 141.665 ;
        RECT 2372.730 131.565 2842.270 135.815 ;
        RECT 2372.730 105.015 2375.000 129.965 ;
      LAYER met5 ;
        RECT 2376.600 105.015 2391.400 129.965 ;
      LAYER met5 ;
        RECT 2393.000 105.015 2395.000 129.965 ;
      LAYER met5 ;
        RECT 2396.600 105.015 2411.400 129.965 ;
      LAYER met5 ;
        RECT 2413.000 105.015 2415.000 129.965 ;
      LAYER met5 ;
        RECT 2416.600 105.015 2431.400 129.965 ;
      LAYER met5 ;
        RECT 2433.000 105.015 2435.000 129.965 ;
      LAYER met5 ;
        RECT 2436.600 105.015 2451.400 129.965 ;
      LAYER met5 ;
        RECT 2453.000 105.015 2455.000 129.965 ;
      LAYER met5 ;
        RECT 2456.600 105.015 2471.400 129.965 ;
      LAYER met5 ;
        RECT 2473.000 105.015 2475.000 129.965 ;
      LAYER met5 ;
        RECT 2476.600 105.015 2491.400 129.965 ;
      LAYER met5 ;
        RECT 2493.000 105.015 2495.000 129.965 ;
      LAYER met5 ;
        RECT 2496.600 105.015 2511.400 129.965 ;
      LAYER met5 ;
        RECT 2513.000 105.015 2515.000 129.965 ;
      LAYER met5 ;
        RECT 2516.600 105.015 2531.400 129.965 ;
      LAYER met5 ;
        RECT 2533.000 105.015 2535.000 129.965 ;
      LAYER met5 ;
        RECT 2536.600 105.015 2551.400 129.965 ;
      LAYER met5 ;
        RECT 2553.000 105.015 2555.000 129.965 ;
      LAYER met5 ;
        RECT 2556.600 105.015 2571.400 129.965 ;
      LAYER met5 ;
        RECT 2573.000 105.015 2575.000 129.965 ;
      LAYER met5 ;
        RECT 2576.600 105.015 2591.400 129.965 ;
      LAYER met5 ;
        RECT 2593.000 105.015 2595.000 129.965 ;
      LAYER met5 ;
        RECT 2596.600 105.015 2611.400 129.965 ;
      LAYER met5 ;
        RECT 2613.000 105.015 2615.000 129.965 ;
      LAYER met5 ;
        RECT 2616.600 105.015 2631.400 129.965 ;
      LAYER met5 ;
        RECT 2633.000 105.015 2635.000 129.965 ;
      LAYER met5 ;
        RECT 2636.600 105.015 2651.400 129.965 ;
      LAYER met5 ;
        RECT 2653.000 105.015 2655.000 129.965 ;
      LAYER met5 ;
        RECT 2656.600 105.015 2671.400 129.965 ;
      LAYER met5 ;
        RECT 2673.000 105.015 2675.000 129.965 ;
      LAYER met5 ;
        RECT 2676.600 105.015 2691.400 129.965 ;
      LAYER met5 ;
        RECT 2693.000 105.015 2695.000 129.965 ;
      LAYER met5 ;
        RECT 2696.600 105.015 2711.400 129.965 ;
      LAYER met5 ;
        RECT 2713.000 105.015 2715.000 129.965 ;
      LAYER met5 ;
        RECT 2716.600 105.015 2731.400 129.965 ;
      LAYER met5 ;
        RECT 2733.000 105.015 2735.000 129.965 ;
      LAYER met5 ;
        RECT 2736.600 105.015 2751.400 129.965 ;
      LAYER met5 ;
        RECT 2753.000 105.015 2755.000 129.965 ;
      LAYER met5 ;
        RECT 2756.600 105.015 2771.400 129.965 ;
      LAYER met5 ;
        RECT 2773.000 105.015 2775.000 129.965 ;
      LAYER met5 ;
        RECT 2776.600 105.015 2791.400 129.965 ;
      LAYER met5 ;
        RECT 2793.000 105.015 2795.000 129.965 ;
      LAYER met5 ;
        RECT 2796.600 105.015 2811.400 129.965 ;
      LAYER met5 ;
        RECT 2813.000 105.015 2815.000 129.965 ;
      LAYER met5 ;
        RECT 2816.600 105.015 2831.400 129.965 ;
      LAYER met5 ;
        RECT 2833.000 105.015 2835.000 129.965 ;
        RECT 2838.000 105.015 2842.270 129.965 ;
      LAYER met5 ;
        RECT 2843.870 103.415 2913.130 181.715 ;
      LAYER met5 ;
        RECT 2914.730 175.665 3385.270 180.115 ;
      LAYER met5 ;
        RECT 3386.870 175.245 3434.135 181.715 ;
      LAYER met5 ;
        RECT 3435.735 176.845 3444.735 729.270 ;
        RECT 3446.335 198.375 3450.585 729.270 ;
        RECT 3452.185 198.520 3456.435 729.270 ;
        RECT 3458.035 724.000 3482.985 729.270 ;
      LAYER met5 ;
        RECT 3484.585 728.000 3588.000 730.870 ;
      LAYER met5 ;
        RECT 3458.035 719.000 3482.985 721.000 ;
      LAYER met5 ;
        RECT 3458.035 702.600 3482.985 717.400 ;
      LAYER met5 ;
        RECT 3458.035 699.000 3482.985 701.000 ;
      LAYER met5 ;
        RECT 3458.035 682.600 3482.985 697.400 ;
      LAYER met5 ;
        RECT 3458.035 679.000 3482.985 681.000 ;
      LAYER met5 ;
        RECT 3458.035 662.600 3482.985 677.400 ;
      LAYER met5 ;
        RECT 3458.035 659.000 3482.985 661.000 ;
      LAYER met5 ;
        RECT 3458.035 642.600 3482.985 657.400 ;
      LAYER met5 ;
        RECT 3458.035 639.000 3482.985 641.000 ;
      LAYER met5 ;
        RECT 3458.035 622.600 3482.985 637.400 ;
      LAYER met5 ;
        RECT 3458.035 619.000 3482.985 621.000 ;
      LAYER met5 ;
        RECT 3458.035 602.600 3482.985 617.400 ;
      LAYER met5 ;
        RECT 3458.035 599.000 3482.985 601.000 ;
      LAYER met5 ;
        RECT 3458.035 582.600 3482.985 597.400 ;
      LAYER met5 ;
        RECT 3458.035 579.000 3482.985 581.000 ;
      LAYER met5 ;
        RECT 3458.035 562.600 3482.985 577.400 ;
      LAYER met5 ;
        RECT 3458.035 559.000 3482.985 561.000 ;
      LAYER met5 ;
        RECT 3458.035 542.600 3482.985 557.400 ;
      LAYER met5 ;
        RECT 3458.035 539.000 3482.985 541.000 ;
      LAYER met5 ;
        RECT 3458.035 522.600 3482.985 537.400 ;
      LAYER met5 ;
        RECT 3458.035 519.000 3482.985 521.000 ;
      LAYER met5 ;
        RECT 3458.035 502.600 3482.985 517.400 ;
      LAYER met5 ;
        RECT 3458.035 499.000 3482.985 501.000 ;
      LAYER met5 ;
        RECT 3458.035 482.600 3482.985 497.400 ;
      LAYER met5 ;
        RECT 3458.035 479.000 3482.985 481.000 ;
      LAYER met5 ;
        RECT 3458.035 462.600 3482.985 477.400 ;
      LAYER met5 ;
        RECT 3458.035 459.000 3482.985 461.000 ;
      LAYER met5 ;
        RECT 3458.035 442.600 3482.985 457.400 ;
      LAYER met5 ;
        RECT 3458.035 439.000 3482.985 441.000 ;
      LAYER met5 ;
        RECT 3458.035 422.600 3482.985 437.400 ;
      LAYER met5 ;
        RECT 3458.035 419.000 3482.985 421.000 ;
      LAYER met5 ;
        RECT 3458.035 402.600 3482.985 417.400 ;
      LAYER met5 ;
        RECT 3458.035 399.000 3482.985 401.000 ;
      LAYER met5 ;
        RECT 3458.035 382.600 3482.985 397.400 ;
      LAYER met5 ;
        RECT 3458.035 379.000 3482.985 381.000 ;
      LAYER met5 ;
        RECT 3458.035 362.600 3482.985 377.400 ;
      LAYER met5 ;
        RECT 3458.035 359.000 3482.985 361.000 ;
      LAYER met5 ;
        RECT 3458.035 342.600 3482.985 357.400 ;
      LAYER met5 ;
        RECT 3458.035 339.000 3482.985 341.000 ;
      LAYER met5 ;
        RECT 3458.035 322.600 3482.985 337.400 ;
      LAYER met5 ;
        RECT 3458.035 319.000 3482.985 321.000 ;
      LAYER met5 ;
        RECT 3458.035 302.600 3482.985 317.400 ;
      LAYER met5 ;
        RECT 3458.035 299.000 3482.985 301.000 ;
      LAYER met5 ;
        RECT 3458.035 282.600 3482.985 297.400 ;
      LAYER met5 ;
        RECT 3458.035 279.000 3482.985 281.000 ;
      LAYER met5 ;
        RECT 3458.035 262.600 3482.985 277.400 ;
      LAYER met5 ;
        RECT 3458.035 259.000 3482.985 261.000 ;
      LAYER met5 ;
        RECT 3458.035 242.600 3482.985 257.400 ;
      LAYER met5 ;
        RECT 3458.035 239.000 3482.985 241.000 ;
      LAYER met5 ;
        RECT 3458.035 222.600 3482.985 237.400 ;
      LAYER met5 ;
        RECT 3458.035 219.000 3482.985 221.000 ;
      LAYER met5 ;
        RECT 3458.035 202.600 3482.985 217.400 ;
      LAYER met5 ;
        RECT 3458.035 197.355 3482.985 201.000 ;
        RECT 3563.785 200.000 3588.000 728.000 ;
      LAYER met5 ;
        RECT 3452.185 196.775 3456.435 196.920 ;
        RECT 3446.335 195.755 3456.435 196.775 ;
        RECT 3484.585 195.755 3588.000 200.000 ;
        RECT 3446.335 175.245 3588.000 195.755 ;
      LAYER met5 ;
        RECT 2914.730 169.615 3385.270 174.065 ;
        RECT 2914.730 164.765 3385.270 168.015 ;
        RECT 2916.000 163.160 3384.000 163.165 ;
        RECT 2914.730 159.915 3385.270 163.160 ;
        RECT 2914.730 153.865 3385.270 158.315 ;
      LAYER met5 ;
        RECT 3386.870 153.865 3588.000 175.245 ;
      LAYER met5 ;
        RECT 2914.730 143.265 3411.155 152.265 ;
      LAYER met5 ;
        RECT 3412.755 141.665 3588.000 153.865 ;
      LAYER met5 ;
        RECT 2914.730 137.415 3385.270 141.665 ;
        RECT 2914.730 131.565 3385.270 135.815 ;
      LAYER met5 ;
        RECT 3386.870 131.565 3588.000 141.665 ;
      LAYER met5 ;
        RECT 2914.730 105.015 2917.000 129.965 ;
      LAYER met5 ;
        RECT 2918.600 105.015 2933.400 129.965 ;
      LAYER met5 ;
        RECT 2935.000 105.015 2937.000 129.965 ;
      LAYER met5 ;
        RECT 2938.600 105.015 2953.400 129.965 ;
      LAYER met5 ;
        RECT 2955.000 105.015 2957.000 129.965 ;
      LAYER met5 ;
        RECT 2958.600 105.015 2973.400 129.965 ;
      LAYER met5 ;
        RECT 2975.000 105.015 2977.000 129.965 ;
      LAYER met5 ;
        RECT 2978.600 105.015 2993.400 129.965 ;
      LAYER met5 ;
        RECT 2995.000 105.015 2997.000 129.965 ;
      LAYER met5 ;
        RECT 2998.600 105.015 3013.400 129.965 ;
      LAYER met5 ;
        RECT 3015.000 105.015 3017.000 129.965 ;
      LAYER met5 ;
        RECT 3018.600 105.015 3033.400 129.965 ;
      LAYER met5 ;
        RECT 3035.000 105.015 3037.000 129.965 ;
      LAYER met5 ;
        RECT 3038.600 105.015 3053.400 129.965 ;
      LAYER met5 ;
        RECT 3055.000 105.015 3057.000 129.965 ;
      LAYER met5 ;
        RECT 3058.600 105.015 3073.400 129.965 ;
      LAYER met5 ;
        RECT 3075.000 105.015 3077.000 129.965 ;
      LAYER met5 ;
        RECT 3078.600 105.015 3093.400 129.965 ;
      LAYER met5 ;
        RECT 3095.000 105.015 3097.000 129.965 ;
      LAYER met5 ;
        RECT 3098.600 105.015 3113.400 129.965 ;
      LAYER met5 ;
        RECT 3115.000 105.015 3117.000 129.965 ;
      LAYER met5 ;
        RECT 3118.600 105.015 3133.400 129.965 ;
      LAYER met5 ;
        RECT 3135.000 105.015 3137.000 129.965 ;
      LAYER met5 ;
        RECT 3138.600 105.015 3153.400 129.965 ;
      LAYER met5 ;
        RECT 3155.000 105.015 3157.000 129.965 ;
      LAYER met5 ;
        RECT 3158.600 105.015 3173.400 129.965 ;
      LAYER met5 ;
        RECT 3175.000 105.015 3177.000 129.965 ;
      LAYER met5 ;
        RECT 3178.600 105.015 3193.400 129.965 ;
      LAYER met5 ;
        RECT 3195.000 105.015 3197.000 129.965 ;
      LAYER met5 ;
        RECT 3198.600 105.015 3213.400 129.965 ;
      LAYER met5 ;
        RECT 3215.000 105.015 3217.000 129.965 ;
      LAYER met5 ;
        RECT 3218.600 105.015 3233.400 129.965 ;
      LAYER met5 ;
        RECT 3235.000 105.015 3237.000 129.965 ;
      LAYER met5 ;
        RECT 3238.600 105.015 3253.400 129.965 ;
      LAYER met5 ;
        RECT 3255.000 105.015 3257.000 129.965 ;
      LAYER met5 ;
        RECT 3258.600 105.015 3273.400 129.965 ;
      LAYER met5 ;
        RECT 3275.000 105.015 3277.000 129.965 ;
      LAYER met5 ;
        RECT 3278.600 105.015 3293.400 129.965 ;
      LAYER met5 ;
        RECT 3295.000 105.015 3297.000 129.965 ;
      LAYER met5 ;
        RECT 3298.600 105.015 3313.400 129.965 ;
      LAYER met5 ;
        RECT 3315.000 105.015 3317.000 129.965 ;
      LAYER met5 ;
        RECT 3318.600 105.015 3333.400 129.965 ;
      LAYER met5 ;
        RECT 3335.000 105.015 3337.000 129.965 ;
      LAYER met5 ;
        RECT 3338.600 105.015 3353.400 129.965 ;
      LAYER met5 ;
        RECT 3355.000 105.015 3357.000 129.965 ;
      LAYER met5 ;
        RECT 3358.600 105.015 3373.400 129.965 ;
      LAYER met5 ;
        RECT 3375.000 105.015 3377.000 129.965 ;
        RECT 3380.000 105.015 3385.855 129.965 ;
      LAYER met5 ;
        RECT 3387.455 103.415 3588.000 131.565 ;
        RECT 0.000 0.000 200.000 103.415 ;
        RECT 667.000 97.590 742.000 103.415 ;
        RECT 667.000 31.775 671.600 97.590 ;
        RECT 737.500 31.775 742.000 97.590 ;
      LAYER met5 ;
        RECT 200.000 0.000 667.000 24.215 ;
      LAYER met5 ;
        RECT 667.000 0.000 742.000 31.775 ;
        RECT 1209.000 97.590 1284.000 103.415 ;
        RECT 1209.000 31.775 1213.600 97.590 ;
        RECT 1279.500 31.775 1284.000 97.590 ;
      LAYER met5 ;
        RECT 742.000 0.000 1209.000 24.215 ;
      LAYER met5 ;
        RECT 1209.000 0.000 1284.000 31.775 ;
        RECT 1752.000 97.040 1832.000 103.415 ;
        RECT 1752.000 31.390 1756.600 97.040 ;
        RECT 1822.400 31.390 1832.000 97.040 ;
      LAYER met5 ;
        RECT 1284.000 0.000 1752.000 24.215 ;
      LAYER met5 ;
        RECT 1752.000 0.000 1832.000 31.390 ;
        RECT 2299.000 99.460 2374.000 103.415 ;
        RECT 2299.000 28.830 2306.445 99.460 ;
        RECT 2366.285 28.830 2374.000 99.460 ;
      LAYER met5 ;
        RECT 1832.000 0.000 2299.000 24.215 ;
      LAYER met5 ;
        RECT 2299.000 0.000 2374.000 28.830 ;
        RECT 2841.000 97.590 2916.000 103.415 ;
        RECT 2841.000 31.775 2845.600 97.590 ;
        RECT 2911.500 31.775 2916.000 97.590 ;
      LAYER met5 ;
        RECT 2374.000 0.000 2841.000 24.215 ;
      LAYER met5 ;
        RECT 2841.000 0.000 2916.000 31.775 ;
      LAYER met5 ;
        RECT 2916.000 0.000 3384.000 24.215 ;
      LAYER met5 ;
        RECT 3384.000 0.000 3588.000 103.415 ;
  END
END chip_io
END LIBRARY

