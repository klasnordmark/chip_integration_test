VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO testdesign
  CLASS BLOCK ;
  FOREIGN testdesign ;
  ORIGIN 0.000 0.000 ;
  SIZE 116.660 BY 115.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 56.345 52.825 56.660 53.385 ;
      LAYER mcon ;
        RECT 56.405 53.165 56.575 53.335 ;
      LAYER met1 ;
        RECT 56.345 53.320 56.635 53.365 ;
        RECT 73.350 53.320 73.670 53.380 ;
        RECT 56.345 53.180 73.670 53.320 ;
        RECT 56.345 53.135 56.635 53.180 ;
        RECT 73.350 53.120 73.670 53.180 ;
      LAYER via ;
        RECT 73.380 53.120 73.640 53.380 ;
      LAYER met2 ;
        RECT 75.670 107.135 75.950 111.135 ;
        RECT 75.740 106.870 75.880 107.135 ;
        RECT 73.440 106.730 75.880 106.870 ;
        RECT 73.440 53.410 73.580 106.730 ;
        RECT 73.380 53.090 73.640 53.410 ;
    END
  END clk
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 60.545 18.095 60.920 18.425 ;
      LAYER mcon ;
        RECT 60.545 18.145 60.715 18.315 ;
      LAYER met1 ;
        RECT 60.485 18.300 60.775 18.345 ;
        RECT 68.290 18.300 68.610 18.360 ;
        RECT 60.485 18.160 68.610 18.300 ;
        RECT 60.485 18.115 60.775 18.160 ;
        RECT 68.290 18.100 68.610 18.160 ;
      LAYER via ;
        RECT 68.320 18.100 68.580 18.360 ;
      LAYER met2 ;
        RECT 68.320 18.070 68.580 18.390 ;
        RECT 68.380 9.820 68.520 18.070 ;
        RECT 68.310 5.820 68.590 9.820 ;
    END
  END in[0]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 60.085 45.295 60.460 45.625 ;
      LAYER mcon ;
        RECT 60.085 45.345 60.255 45.515 ;
      LAYER met1 ;
        RECT 60.010 45.500 60.330 45.560 ;
        RECT 59.815 45.360 60.330 45.500 ;
        RECT 60.010 45.300 60.330 45.360 ;
        RECT 22.290 23.060 22.610 23.120 ;
        RECT 60.010 23.060 60.330 23.120 ;
        RECT 22.290 22.920 60.330 23.060 ;
        RECT 22.290 22.860 22.610 22.920 ;
        RECT 60.010 22.860 60.330 22.920 ;
      LAYER via ;
        RECT 60.040 45.300 60.300 45.560 ;
        RECT 22.320 22.860 22.580 23.120 ;
        RECT 60.040 22.860 60.300 23.120 ;
      LAYER met2 ;
        RECT 60.040 45.270 60.300 45.590 ;
        RECT 60.100 23.150 60.240 45.270 ;
        RECT 22.320 22.830 22.580 23.150 ;
        RECT 60.040 22.830 60.300 23.150 ;
        RECT 22.380 9.820 22.520 22.830 ;
        RECT 22.310 5.820 22.590 9.820 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 65.605 56.175 65.980 56.505 ;
      LAYER mcon ;
        RECT 65.605 56.225 65.775 56.395 ;
      LAYER met1 ;
        RECT 17.690 56.380 18.010 56.440 ;
        RECT 65.545 56.380 65.835 56.425 ;
        RECT 17.690 56.240 65.835 56.380 ;
        RECT 17.690 56.180 18.010 56.240 ;
        RECT 65.545 56.195 65.835 56.240 ;
        RECT 14.010 23.400 14.330 23.460 ;
        RECT 17.690 23.400 18.010 23.460 ;
        RECT 14.010 23.260 18.010 23.400 ;
        RECT 14.010 23.200 14.330 23.260 ;
        RECT 17.690 23.200 18.010 23.260 ;
      LAYER via ;
        RECT 17.720 56.180 17.980 56.440 ;
        RECT 14.040 23.200 14.300 23.460 ;
        RECT 17.720 23.200 17.980 23.460 ;
      LAYER met2 ;
        RECT 17.720 56.150 17.980 56.470 ;
        RECT 17.780 23.490 17.920 56.150 ;
        RECT 14.040 23.170 14.300 23.490 ;
        RECT 17.720 23.170 17.980 23.490 ;
        RECT 14.100 9.820 14.240 23.170 ;
        RECT 14.030 5.820 14.310 9.820 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 64.685 91.135 65.060 91.465 ;
      LAYER mcon ;
        RECT 64.685 91.245 64.855 91.415 ;
      LAYER met1 ;
        RECT 64.625 91.400 64.915 91.445 ;
        RECT 94.050 91.400 94.370 91.460 ;
        RECT 64.625 91.260 94.370 91.400 ;
        RECT 64.625 91.215 64.915 91.260 ;
        RECT 94.050 91.200 94.370 91.260 ;
      LAYER via ;
        RECT 94.080 91.200 94.340 91.460 ;
      LAYER met2 ;
        RECT 94.070 107.135 94.350 111.135 ;
        RECT 94.140 91.490 94.280 107.135 ;
        RECT 94.080 91.170 94.340 91.490 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 64.225 58.495 64.600 58.825 ;
      LAYER mcon ;
        RECT 64.225 58.605 64.395 58.775 ;
      LAYER met1 ;
        RECT 64.165 58.760 64.455 58.805 ;
        RECT 94.050 58.760 94.370 58.820 ;
        RECT 64.165 58.620 94.370 58.760 ;
        RECT 64.165 58.575 64.455 58.620 ;
        RECT 94.050 58.560 94.370 58.620 ;
      LAYER via ;
        RECT 94.080 58.560 94.340 58.820 ;
      LAYER met2 ;
        RECT 94.080 58.530 94.340 58.850 ;
        RECT 94.140 10.310 94.280 58.530 ;
        RECT 94.140 10.170 95.200 10.310 ;
        RECT 95.060 9.820 95.200 10.170 ;
        RECT 94.990 5.820 95.270 9.820 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 73.425 23.535 73.800 23.865 ;
      LAYER mcon ;
        RECT 73.425 23.585 73.595 23.755 ;
      LAYER met1 ;
        RECT 73.365 23.740 73.655 23.785 ;
        RECT 80.250 23.740 80.570 23.800 ;
        RECT 73.365 23.600 80.570 23.740 ;
        RECT 73.365 23.555 73.655 23.600 ;
        RECT 80.250 23.540 80.570 23.600 ;
      LAYER via ;
        RECT 80.280 23.540 80.540 23.800 ;
      LAYER met2 ;
        RECT 80.270 25.015 80.550 25.385 ;
        RECT 80.340 23.830 80.480 25.015 ;
        RECT 80.280 23.510 80.540 23.830 ;
      LAYER via2 ;
        RECT 80.270 25.060 80.550 25.340 ;
      LAYER met3 ;
        RECT 80.245 25.350 80.575 25.365 ;
        RECT 101.775 25.350 105.775 25.500 ;
        RECT 80.245 25.050 105.775 25.350 ;
        RECT 80.245 25.035 80.575 25.050 ;
        RECT 101.775 24.900 105.775 25.050 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 37.985 58.495 38.295 59.115 ;
      LAYER mcon ;
        RECT 38.005 58.605 38.175 58.775 ;
      LAYER met1 ;
        RECT 37.945 58.760 38.235 58.805 ;
        RECT 37.560 58.620 38.235 58.760 ;
        RECT 37.560 58.080 37.700 58.620 ;
        RECT 37.945 58.575 38.235 58.620 ;
        RECT 38.850 58.080 39.170 58.140 ;
        RECT 37.560 57.940 39.170 58.080 ;
        RECT 38.850 57.880 39.170 57.940 ;
      LAYER via ;
        RECT 38.880 57.880 39.140 58.140 ;
      LAYER met2 ;
        RECT 38.880 57.850 39.140 58.170 ;
        RECT 38.940 10.310 39.080 57.850 ;
        RECT 38.940 10.170 40.920 10.310 ;
        RECT 40.780 9.820 40.920 10.170 ;
        RECT 40.710 5.820 40.990 9.820 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 38.465 80.255 38.840 80.585 ;
      LAYER mcon ;
        RECT 38.465 80.365 38.635 80.535 ;
      LAYER met1 ;
        RECT 38.390 80.520 38.710 80.580 ;
        RECT 38.390 80.380 38.905 80.520 ;
        RECT 38.390 80.320 38.710 80.380 ;
      LAYER via ;
        RECT 38.420 80.320 38.680 80.580 ;
      LAYER met2 ;
        RECT 38.870 107.135 39.150 111.135 ;
        RECT 38.940 106.870 39.080 107.135 ;
        RECT 38.940 106.730 39.540 106.870 ;
        RECT 39.400 95.310 39.540 106.730 ;
        RECT 38.480 95.170 39.540 95.310 ;
        RECT 38.480 80.610 38.620 95.170 ;
        RECT 38.420 80.290 38.680 80.610 ;
    END
  END in[7]
  PIN oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.235 93.115 20.755 94.665 ;
      LAYER mcon ;
        RECT 20.525 94.305 20.695 94.475 ;
      LAYER met1 ;
        RECT 20.465 94.460 20.755 94.505 ;
        RECT 25.050 94.460 25.370 94.520 ;
        RECT 20.465 94.320 25.370 94.460 ;
        RECT 20.465 94.275 20.755 94.320 ;
        RECT 25.050 94.260 25.370 94.320 ;
      LAYER via ;
        RECT 25.080 94.260 25.340 94.520 ;
      LAYER met2 ;
        RECT 25.070 103.895 25.350 104.265 ;
        RECT 25.140 94.550 25.280 103.895 ;
        RECT 25.080 94.230 25.340 94.550 ;
      LAYER via2 ;
        RECT 25.070 103.940 25.350 104.220 ;
      LAYER met3 ;
        RECT 11.180 104.230 15.180 104.380 ;
        RECT 25.045 104.230 25.375 104.245 ;
        RECT 11.180 103.930 25.375 104.230 ;
        RECT 11.180 103.780 15.180 103.930 ;
        RECT 25.045 103.915 25.375 103.930 ;
    END
  END oeb[0]
  PIN oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 60.255 93.115 60.775 94.665 ;
      LAYER mcon ;
        RECT 60.545 94.305 60.715 94.475 ;
      LAYER met1 ;
        RECT 56.790 94.460 57.110 94.520 ;
        RECT 60.485 94.460 60.775 94.505 ;
        RECT 56.790 94.320 60.775 94.460 ;
        RECT 56.790 94.260 57.110 94.320 ;
        RECT 60.485 94.275 60.775 94.320 ;
      LAYER via ;
        RECT 56.820 94.260 57.080 94.520 ;
      LAYER met2 ;
        RECT 57.270 107.135 57.550 111.135 ;
        RECT 57.340 99.390 57.480 107.135 ;
        RECT 56.880 99.250 57.480 99.390 ;
        RECT 56.880 94.550 57.020 99.250 ;
        RECT 56.820 94.230 57.080 94.550 ;
    END
  END oeb[10]
  PIN oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.235 33.275 20.755 34.825 ;
      LAYER mcon ;
        RECT 20.525 34.465 20.695 34.635 ;
      LAYER met1 ;
        RECT 20.450 34.620 20.770 34.680 ;
        RECT 20.255 34.480 20.770 34.620 ;
        RECT 20.450 34.420 20.770 34.480 ;
      LAYER via ;
        RECT 20.480 34.420 20.740 34.680 ;
      LAYER met2 ;
        RECT 20.470 35.895 20.750 36.265 ;
        RECT 20.540 34.710 20.680 35.895 ;
        RECT 20.480 34.390 20.740 34.710 ;
      LAYER via2 ;
        RECT 20.470 35.940 20.750 36.220 ;
      LAYER met3 ;
        RECT 11.180 36.230 15.180 36.380 ;
        RECT 20.445 36.230 20.775 36.245 ;
        RECT 11.180 35.930 20.775 36.230 ;
        RECT 11.180 35.780 15.180 35.930 ;
        RECT 20.445 35.915 20.775 35.930 ;
    END
  END oeb[11]
  PIN oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 94.295 36.655 94.815 38.205 ;
      LAYER mcon ;
        RECT 94.585 37.865 94.755 38.035 ;
      LAYER met1 ;
        RECT 94.510 38.020 94.830 38.080 ;
        RECT 94.315 37.880 94.830 38.020 ;
        RECT 94.510 37.820 94.830 37.880 ;
      LAYER via ;
        RECT 94.540 37.820 94.800 38.080 ;
      LAYER met2 ;
        RECT 94.530 38.615 94.810 38.985 ;
        RECT 94.600 38.110 94.740 38.615 ;
        RECT 94.540 37.790 94.800 38.110 ;
      LAYER via2 ;
        RECT 94.530 38.660 94.810 38.940 ;
      LAYER met3 ;
        RECT 94.505 38.950 94.835 38.965 ;
        RECT 101.775 38.950 105.775 39.100 ;
        RECT 94.505 38.650 105.775 38.950 ;
        RECT 94.505 38.635 94.835 38.650 ;
        RECT 101.775 38.500 105.775 38.650 ;
    END
  END oeb[12]
  PIN oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 94.295 16.955 94.815 18.505 ;
      LAYER mcon ;
        RECT 94.585 17.125 94.755 17.295 ;
      LAYER met1 ;
        RECT 93.590 17.280 93.910 17.340 ;
        RECT 94.525 17.280 94.815 17.325 ;
        RECT 93.590 17.140 94.815 17.280 ;
        RECT 93.590 17.080 93.910 17.140 ;
        RECT 94.525 17.095 94.815 17.140 ;
      LAYER via ;
        RECT 93.620 17.080 93.880 17.340 ;
      LAYER met2 ;
        RECT 93.620 17.050 93.880 17.370 ;
        RECT 93.680 11.785 93.820 17.050 ;
        RECT 93.610 11.415 93.890 11.785 ;
      LAYER via2 ;
        RECT 93.610 11.460 93.890 11.740 ;
      LAYER met3 ;
        RECT 93.585 11.750 93.915 11.765 ;
        RECT 101.775 11.750 105.775 11.900 ;
        RECT 93.585 11.450 105.775 11.750 ;
        RECT 93.585 11.435 93.915 11.450 ;
        RECT 101.775 11.300 105.775 11.450 ;
    END
  END oeb[13]
  PIN oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.235 20.335 20.755 21.885 ;
      LAYER mcon ;
        RECT 20.525 21.545 20.695 21.715 ;
      LAYER met1 ;
        RECT 20.450 21.700 20.770 21.760 ;
        RECT 20.255 21.560 20.770 21.700 ;
        RECT 20.450 21.500 20.770 21.560 ;
      LAYER via ;
        RECT 20.480 21.500 20.740 21.760 ;
      LAYER met2 ;
        RECT 20.470 22.295 20.750 22.665 ;
        RECT 20.540 21.790 20.680 22.295 ;
        RECT 20.480 21.470 20.740 21.790 ;
      LAYER via2 ;
        RECT 20.470 22.340 20.750 22.620 ;
      LAYER met3 ;
        RECT 11.180 22.630 15.180 22.780 ;
        RECT 20.445 22.630 20.775 22.645 ;
        RECT 11.180 22.330 20.775 22.630 ;
        RECT 11.180 22.180 15.180 22.330 ;
        RECT 20.445 22.315 20.775 22.330 ;
    END
  END oeb[14]
  PIN oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 32.195 16.955 32.715 18.505 ;
      LAYER mcon ;
        RECT 32.485 17.125 32.655 17.295 ;
      LAYER met1 ;
        RECT 31.490 17.280 31.810 17.340 ;
        RECT 32.425 17.280 32.715 17.325 ;
        RECT 31.490 17.140 32.715 17.280 ;
        RECT 31.490 17.080 31.810 17.140 ;
        RECT 32.425 17.095 32.715 17.140 ;
      LAYER via ;
        RECT 31.520 17.080 31.780 17.340 ;
      LAYER met2 ;
        RECT 31.520 17.050 31.780 17.370 ;
        RECT 31.580 9.820 31.720 17.050 ;
        RECT 31.510 5.820 31.790 9.820 ;
    END
  END oeb[15]
  PIN oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 94.295 93.115 94.815 94.665 ;
      LAYER mcon ;
        RECT 94.585 94.305 94.755 94.475 ;
      LAYER met1 ;
        RECT 94.525 94.460 94.815 94.505 ;
        RECT 102.330 94.460 102.650 94.520 ;
        RECT 94.525 94.320 102.650 94.460 ;
        RECT 94.525 94.275 94.815 94.320 ;
        RECT 102.330 94.260 102.650 94.320 ;
      LAYER via ;
        RECT 102.360 94.260 102.620 94.520 ;
      LAYER met2 ;
        RECT 102.350 107.135 102.630 111.135 ;
        RECT 102.420 94.550 102.560 107.135 ;
        RECT 102.360 94.230 102.620 94.550 ;
    END
  END oeb[1]
  PIN oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.235 47.535 20.755 49.085 ;
      LAYER mcon ;
        RECT 20.525 48.745 20.695 48.915 ;
      LAYER met1 ;
        RECT 20.450 48.900 20.770 48.960 ;
        RECT 20.255 48.760 20.770 48.900 ;
        RECT 20.450 48.700 20.770 48.760 ;
      LAYER via ;
        RECT 20.480 48.700 20.740 48.960 ;
      LAYER met2 ;
        RECT 20.470 49.495 20.750 49.865 ;
        RECT 20.540 48.990 20.680 49.495 ;
        RECT 20.480 48.670 20.740 48.990 ;
      LAYER via2 ;
        RECT 20.470 49.540 20.750 49.820 ;
      LAYER met3 ;
        RECT 11.180 49.830 15.180 49.980 ;
        RECT 20.445 49.830 20.775 49.845 ;
        RECT 11.180 49.530 20.775 49.830 ;
        RECT 11.180 49.380 15.180 49.530 ;
        RECT 20.445 49.515 20.775 49.530 ;
    END
  END oeb[2]
  PIN oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 88.315 93.115 88.835 94.665 ;
      LAYER mcon ;
        RECT 88.605 94.305 88.775 94.475 ;
      LAYER met1 ;
        RECT 84.850 94.460 85.170 94.520 ;
        RECT 88.545 94.460 88.835 94.505 ;
        RECT 84.850 94.320 88.835 94.460 ;
        RECT 84.850 94.260 85.170 94.320 ;
        RECT 88.545 94.275 88.835 94.320 ;
      LAYER via ;
        RECT 84.880 94.260 85.140 94.520 ;
      LAYER met2 ;
        RECT 84.870 107.135 85.150 111.135 ;
        RECT 84.940 94.550 85.080 107.135 ;
        RECT 84.880 94.230 85.140 94.550 ;
    END
  END oeb[3]
  PIN oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 32.195 93.115 32.715 94.665 ;
      LAYER mcon ;
        RECT 32.485 94.305 32.655 94.475 ;
      LAYER met1 ;
        RECT 29.190 94.460 29.510 94.520 ;
        RECT 32.425 94.460 32.715 94.505 ;
        RECT 29.190 94.320 32.715 94.460 ;
        RECT 29.190 94.260 29.510 94.320 ;
        RECT 32.425 94.275 32.715 94.320 ;
      LAYER via ;
        RECT 29.220 94.260 29.480 94.520 ;
      LAYER met2 ;
        RECT 29.670 107.135 29.950 111.135 ;
        RECT 29.740 99.390 29.880 107.135 ;
        RECT 29.280 99.250 29.880 99.390 ;
        RECT 29.280 94.550 29.420 99.250 ;
        RECT 29.220 94.230 29.480 94.550 ;
    END
  END oeb[4]
  PIN oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 94.295 91.055 94.815 92.605 ;
      LAYER mcon ;
        RECT 94.585 92.265 94.755 92.435 ;
      LAYER met1 ;
        RECT 94.510 92.420 94.830 92.480 ;
        RECT 94.315 92.280 94.830 92.420 ;
        RECT 94.510 92.220 94.830 92.280 ;
      LAYER via ;
        RECT 94.540 92.220 94.800 92.480 ;
      LAYER met2 ;
        RECT 94.530 93.015 94.810 93.385 ;
        RECT 94.600 92.510 94.740 93.015 ;
        RECT 94.540 92.190 94.800 92.510 ;
      LAYER via2 ;
        RECT 94.530 93.060 94.810 93.340 ;
      LAYER met3 ;
        RECT 94.505 93.350 94.835 93.365 ;
        RECT 101.775 93.350 105.775 93.500 ;
        RECT 94.505 93.050 105.775 93.350 ;
        RECT 94.505 93.035 94.835 93.050 ;
        RECT 101.775 92.900 105.775 93.050 ;
    END
  END oeb[5]
  PIN oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 89.235 16.955 89.755 18.505 ;
      LAYER mcon ;
        RECT 89.525 17.125 89.695 17.295 ;
      LAYER met1 ;
        RECT 87.150 17.280 87.470 17.340 ;
        RECT 89.465 17.280 89.755 17.325 ;
        RECT 87.150 17.140 89.755 17.280 ;
        RECT 87.150 17.080 87.470 17.140 ;
        RECT 89.465 17.095 89.755 17.140 ;
      LAYER via ;
        RECT 87.180 17.080 87.440 17.340 ;
      LAYER met2 ;
        RECT 87.180 17.050 87.440 17.370 ;
        RECT 87.240 13.030 87.380 17.050 ;
        RECT 86.780 12.890 87.380 13.030 ;
        RECT 86.780 9.820 86.920 12.890 ;
        RECT 86.710 5.820 86.990 9.820 ;
    END
  END oeb[6]
  PIN oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.235 60.475 20.755 62.025 ;
      LAYER mcon ;
        RECT 20.525 61.665 20.695 61.835 ;
      LAYER met1 ;
        RECT 20.450 61.820 20.770 61.880 ;
        RECT 20.255 61.680 20.770 61.820 ;
        RECT 20.450 61.620 20.770 61.680 ;
      LAYER via ;
        RECT 20.480 61.620 20.740 61.880 ;
      LAYER met2 ;
        RECT 20.470 63.095 20.750 63.465 ;
        RECT 20.540 61.910 20.680 63.095 ;
        RECT 20.480 61.590 20.740 61.910 ;
      LAYER via2 ;
        RECT 20.470 63.140 20.750 63.420 ;
      LAYER met3 ;
        RECT 11.180 63.430 15.180 63.580 ;
        RECT 20.445 63.430 20.775 63.445 ;
        RECT 11.180 63.130 20.775 63.430 ;
        RECT 11.180 62.980 15.180 63.130 ;
        RECT 20.445 63.115 20.775 63.130 ;
    END
  END oeb[7]
  PIN oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 80.265 78.530 80.600 78.955 ;
        RECT 81.120 78.530 81.455 78.955 ;
        RECT 80.265 78.360 81.935 78.530 ;
        RECT 81.690 77.795 81.935 78.360 ;
        RECT 80.265 77.625 81.935 77.795 ;
        RECT 80.265 76.865 80.600 77.625 ;
        RECT 81.120 76.865 81.450 77.625 ;
      LAYER mcon ;
        RECT 81.705 78.325 81.875 78.495 ;
      LAYER met1 ;
        RECT 81.630 78.480 81.950 78.540 ;
        RECT 81.435 78.340 81.950 78.480 ;
        RECT 81.630 78.280 81.950 78.340 ;
      LAYER via ;
        RECT 81.660 78.280 81.920 78.540 ;
      LAYER met2 ;
        RECT 81.650 79.415 81.930 79.785 ;
        RECT 81.720 78.570 81.860 79.415 ;
        RECT 81.660 78.250 81.920 78.570 ;
      LAYER via2 ;
        RECT 81.650 79.460 81.930 79.740 ;
      LAYER met3 ;
        RECT 81.625 79.750 81.955 79.765 ;
        RECT 101.775 79.750 105.775 79.900 ;
        RECT 81.625 79.450 105.775 79.750 ;
        RECT 81.625 79.435 81.955 79.450 ;
        RECT 101.775 79.300 105.775 79.450 ;
    END
  END oeb[8]
  PIN oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 49.675 16.955 50.195 18.505 ;
      LAYER mcon ;
        RECT 49.965 17.125 50.135 17.295 ;
      LAYER met1 ;
        RECT 49.890 17.280 50.210 17.340 ;
        RECT 49.695 17.140 50.210 17.280 ;
        RECT 49.890 17.080 50.210 17.140 ;
      LAYER via ;
        RECT 49.920 17.080 50.180 17.340 ;
      LAYER met2 ;
        RECT 49.920 17.050 50.180 17.370 ;
        RECT 49.980 9.820 50.120 17.050 ;
        RECT 49.910 5.820 50.190 9.820 ;
    END
  END oeb[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 60.945 21.055 61.280 21.815 ;
        RECT 61.800 21.055 62.130 21.815 ;
        RECT 60.945 20.885 62.615 21.055 ;
        RECT 62.370 20.320 62.615 20.885 ;
        RECT 60.945 20.150 62.615 20.320 ;
        RECT 60.945 19.725 61.280 20.150 ;
        RECT 61.800 19.725 62.135 20.150 ;
      LAYER mcon ;
        RECT 61.005 19.845 61.175 20.015 ;
      LAYER met1 ;
        RECT 59.090 20.000 59.410 20.060 ;
        RECT 60.945 20.000 61.235 20.045 ;
        RECT 59.090 19.860 61.235 20.000 ;
        RECT 59.090 19.800 59.410 19.860 ;
        RECT 60.945 19.815 61.235 19.860 ;
      LAYER via ;
        RECT 59.120 19.800 59.380 20.060 ;
      LAYER met2 ;
        RECT 59.120 19.770 59.380 20.090 ;
        RECT 59.180 17.790 59.320 19.770 ;
        RECT 59.180 17.650 59.780 17.790 ;
        RECT 59.640 15.750 59.780 17.650 ;
        RECT 59.180 15.610 59.780 15.750 ;
        RECT 59.180 9.820 59.320 15.610 ;
        RECT 59.110 5.820 59.390 9.820 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 67.845 51.330 68.180 51.755 ;
        RECT 68.700 51.330 69.035 51.755 ;
        RECT 67.845 51.160 69.515 51.330 ;
        RECT 69.270 50.595 69.515 51.160 ;
        RECT 67.845 50.425 69.515 50.595 ;
        RECT 67.845 49.665 68.180 50.425 ;
        RECT 68.700 49.665 69.030 50.425 ;
      LAYER mcon ;
        RECT 69.285 51.125 69.455 51.295 ;
      LAYER met1 ;
        RECT 69.225 51.280 69.515 51.325 ;
        RECT 86.690 51.280 87.010 51.340 ;
        RECT 69.225 51.140 87.010 51.280 ;
        RECT 69.225 51.095 69.515 51.140 ;
        RECT 86.690 51.080 87.010 51.140 ;
      LAYER via ;
        RECT 86.720 51.080 86.980 51.340 ;
      LAYER met2 ;
        RECT 86.710 52.215 86.990 52.585 ;
        RECT 86.780 51.370 86.920 52.215 ;
        RECT 86.720 51.050 86.980 51.370 ;
      LAYER via2 ;
        RECT 86.710 52.260 86.990 52.540 ;
      LAYER met3 ;
        RECT 86.685 52.550 87.015 52.565 ;
        RECT 101.775 52.550 105.775 52.700 ;
        RECT 86.685 52.250 105.775 52.550 ;
        RECT 86.685 52.235 87.015 52.250 ;
        RECT 101.775 52.100 105.775 52.250 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 75.665 62.210 76.000 62.635 ;
        RECT 76.520 62.210 76.855 62.635 ;
        RECT 75.665 62.040 77.335 62.210 ;
        RECT 77.090 61.475 77.335 62.040 ;
        RECT 75.665 61.305 77.335 61.475 ;
        RECT 75.665 60.545 76.000 61.305 ;
        RECT 76.520 60.545 76.850 61.305 ;
      LAYER mcon ;
        RECT 77.105 62.005 77.275 62.175 ;
      LAYER met1 ;
        RECT 77.045 62.160 77.335 62.205 ;
        RECT 80.250 62.160 80.570 62.220 ;
        RECT 77.045 62.020 80.570 62.160 ;
        RECT 77.045 61.975 77.335 62.020 ;
        RECT 80.250 61.960 80.570 62.020 ;
      LAYER via ;
        RECT 80.280 61.960 80.540 62.220 ;
      LAYER met2 ;
        RECT 80.270 64.455 80.550 64.825 ;
        RECT 80.340 62.250 80.480 64.455 ;
        RECT 80.280 61.930 80.540 62.250 ;
      LAYER via2 ;
        RECT 80.270 64.500 80.550 64.780 ;
      LAYER met3 ;
        RECT 101.775 66.150 105.775 66.300 ;
        RECT 87.850 65.850 105.775 66.150 ;
        RECT 80.245 64.790 80.575 64.805 ;
        RECT 87.850 64.790 88.150 65.850 ;
        RECT 101.775 65.700 105.775 65.850 ;
        RECT 80.245 64.490 88.150 64.790 ;
        RECT 80.245 64.475 80.575 64.490 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 69.225 89.410 69.560 89.835 ;
        RECT 70.080 89.410 70.415 89.835 ;
        RECT 69.225 89.240 70.895 89.410 ;
        RECT 70.650 88.675 70.895 89.240 ;
        RECT 69.225 88.505 70.895 88.675 ;
        RECT 69.225 87.745 69.560 88.505 ;
        RECT 70.080 87.745 70.410 88.505 ;
      LAYER mcon ;
        RECT 69.285 89.545 69.455 89.715 ;
      LAYER met1 ;
        RECT 28.270 89.700 28.590 89.760 ;
        RECT 69.225 89.700 69.515 89.745 ;
        RECT 28.270 89.560 69.515 89.700 ;
        RECT 28.270 89.500 28.590 89.560 ;
        RECT 69.225 89.515 69.515 89.560 ;
      LAYER via ;
        RECT 28.300 89.500 28.560 89.760 ;
      LAYER met2 ;
        RECT 28.290 90.295 28.570 90.665 ;
        RECT 28.360 89.790 28.500 90.295 ;
        RECT 28.300 89.470 28.560 89.790 ;
      LAYER via2 ;
        RECT 28.290 90.340 28.570 90.620 ;
      LAYER met3 ;
        RECT 11.180 90.630 15.180 90.780 ;
        RECT 28.265 90.630 28.595 90.645 ;
        RECT 11.180 90.330 28.595 90.630 ;
        RECT 11.180 90.180 15.180 90.330 ;
        RECT 28.265 90.315 28.595 90.330 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 67.385 64.575 67.720 65.335 ;
        RECT 68.240 64.575 68.570 65.335 ;
        RECT 67.385 64.405 69.055 64.575 ;
        RECT 68.810 63.840 69.055 64.405 ;
        RECT 67.385 63.670 69.055 63.840 ;
        RECT 67.385 63.245 67.720 63.670 ;
        RECT 68.240 63.245 68.575 63.670 ;
      LAYER mcon ;
        RECT 67.445 65.065 67.615 65.235 ;
      LAYER met1 ;
        RECT 66.450 65.220 66.770 65.280 ;
        RECT 67.385 65.220 67.675 65.265 ;
        RECT 66.450 65.080 67.675 65.220 ;
        RECT 66.450 65.020 66.770 65.080 ;
        RECT 67.385 65.035 67.675 65.080 ;
      LAYER via ;
        RECT 66.480 65.020 66.740 65.280 ;
      LAYER met2 ;
        RECT 66.470 107.135 66.750 111.135 ;
        RECT 66.540 65.310 66.680 107.135 ;
        RECT 66.480 64.990 66.740 65.310 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 80.265 21.055 80.600 21.815 ;
        RECT 81.120 21.055 81.450 21.815 ;
        RECT 80.265 20.885 81.935 21.055 ;
        RECT 81.690 20.320 81.935 20.885 ;
        RECT 80.265 20.150 81.935 20.320 ;
        RECT 80.265 19.725 80.600 20.150 ;
        RECT 81.120 19.725 81.455 20.150 ;
      LAYER mcon ;
        RECT 80.325 19.845 80.495 20.015 ;
      LAYER met1 ;
        RECT 77.950 20.000 78.270 20.060 ;
        RECT 80.265 20.000 80.555 20.045 ;
        RECT 77.950 19.860 80.555 20.000 ;
        RECT 77.950 19.800 78.270 19.860 ;
        RECT 80.265 19.815 80.555 19.860 ;
      LAYER via ;
        RECT 77.980 19.800 78.240 20.060 ;
      LAYER met2 ;
        RECT 77.980 19.770 78.240 20.090 ;
        RECT 78.040 13.030 78.180 19.770 ;
        RECT 77.580 12.890 78.180 13.030 ;
        RECT 77.580 9.820 77.720 12.890 ;
        RECT 77.510 5.820 77.790 9.820 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 47.605 62.210 47.940 62.635 ;
        RECT 48.460 62.210 48.795 62.635 ;
        RECT 47.605 62.040 49.275 62.210 ;
        RECT 49.030 61.475 49.275 62.040 ;
        RECT 47.605 61.305 49.275 61.475 ;
        RECT 47.605 60.545 47.940 61.305 ;
        RECT 48.460 60.545 48.790 61.305 ;
      LAYER mcon ;
        RECT 47.665 62.345 47.835 62.515 ;
      LAYER met1 ;
        RECT 45.750 95.140 46.070 95.200 ;
        RECT 48.050 95.140 48.370 95.200 ;
        RECT 45.750 95.000 48.370 95.140 ;
        RECT 45.750 94.940 46.070 95.000 ;
        RECT 48.050 94.940 48.370 95.000 ;
        RECT 45.750 62.500 46.070 62.560 ;
        RECT 47.605 62.500 47.895 62.545 ;
        RECT 45.750 62.360 47.895 62.500 ;
        RECT 45.750 62.300 46.070 62.360 ;
        RECT 47.605 62.315 47.895 62.360 ;
      LAYER via ;
        RECT 45.780 94.940 46.040 95.200 ;
        RECT 48.080 94.940 48.340 95.200 ;
        RECT 45.780 62.300 46.040 62.560 ;
      LAYER met2 ;
        RECT 48.070 107.135 48.350 111.135 ;
        RECT 48.140 95.230 48.280 107.135 ;
        RECT 45.780 94.910 46.040 95.230 ;
        RECT 48.080 94.910 48.340 95.230 ;
        RECT 45.840 62.590 45.980 94.910 ;
        RECT 45.780 62.270 46.040 62.590 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 45.765 78.530 46.100 78.955 ;
        RECT 46.620 78.530 46.955 78.955 ;
        RECT 45.765 78.360 47.435 78.530 ;
        RECT 47.190 77.795 47.435 78.360 ;
        RECT 45.765 77.625 47.435 77.795 ;
        RECT 45.765 76.865 46.100 77.625 ;
        RECT 46.620 76.865 46.950 77.625 ;
      LAYER mcon ;
        RECT 45.825 76.965 45.995 77.135 ;
      LAYER met1 ;
        RECT 28.270 77.120 28.590 77.180 ;
        RECT 45.765 77.120 46.055 77.165 ;
        RECT 28.270 76.980 46.055 77.120 ;
        RECT 28.270 76.920 28.590 76.980 ;
        RECT 45.765 76.935 46.055 76.980 ;
      LAYER via ;
        RECT 28.300 76.920 28.560 77.180 ;
      LAYER met2 ;
        RECT 28.300 77.065 28.560 77.210 ;
        RECT 28.290 76.695 28.570 77.065 ;
      LAYER via2 ;
        RECT 28.290 76.740 28.570 77.020 ;
      LAYER met3 ;
        RECT 11.180 77.030 15.180 77.180 ;
        RECT 28.265 77.030 28.595 77.045 ;
        RECT 11.180 76.730 28.595 77.030 ;
        RECT 11.180 76.580 15.180 76.730 ;
        RECT 28.265 76.715 28.595 76.730 ;
    END
  END out[7]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 35.205 83.375 35.535 83.625 ;
      LAYER mcon ;
        RECT 35.245 83.425 35.415 83.595 ;
      LAYER met1 ;
        RECT 21.370 91.060 21.690 91.120 ;
        RECT 35.170 91.060 35.490 91.120 ;
        RECT 21.370 90.920 35.490 91.060 ;
        RECT 21.370 90.860 21.690 90.920 ;
        RECT 35.170 90.860 35.490 90.920 ;
        RECT 35.170 83.580 35.490 83.640 ;
        RECT 34.975 83.440 35.490 83.580 ;
        RECT 35.170 83.380 35.490 83.440 ;
      LAYER via ;
        RECT 21.400 90.860 21.660 91.120 ;
        RECT 35.200 90.860 35.460 91.120 ;
        RECT 35.200 83.380 35.460 83.640 ;
      LAYER met2 ;
        RECT 21.390 107.135 21.670 111.135 ;
        RECT 21.460 91.150 21.600 107.135 ;
        RECT 21.400 90.830 21.660 91.150 ;
        RECT 35.200 90.830 35.460 91.150 ;
        RECT 35.260 83.670 35.400 90.830 ;
        RECT 35.200 83.350 35.460 83.670 ;
    END
  END reset
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 16.845 98.215 17.015 98.385 ;
        RECT 17.305 98.215 17.475 98.385 ;
        RECT 17.765 98.215 17.935 98.385 ;
        RECT 18.225 98.215 18.395 98.385 ;
        RECT 18.685 98.215 18.855 98.385 ;
        RECT 19.145 98.215 19.315 98.385 ;
        RECT 19.605 98.215 19.775 98.385 ;
        RECT 20.065 98.215 20.235 98.385 ;
        RECT 20.525 98.215 20.695 98.385 ;
        RECT 20.985 98.215 21.155 98.385 ;
        RECT 21.445 98.215 21.615 98.385 ;
        RECT 21.905 98.215 22.075 98.385 ;
        RECT 22.365 98.215 22.535 98.385 ;
        RECT 22.825 98.215 22.995 98.385 ;
        RECT 23.285 98.215 23.455 98.385 ;
        RECT 23.745 98.215 23.915 98.385 ;
        RECT 24.205 98.215 24.375 98.385 ;
        RECT 24.665 98.215 24.835 98.385 ;
        RECT 25.125 98.215 25.295 98.385 ;
        RECT 25.585 98.215 25.755 98.385 ;
        RECT 26.045 98.215 26.215 98.385 ;
        RECT 26.505 98.215 26.675 98.385 ;
        RECT 26.965 98.215 27.135 98.385 ;
        RECT 27.425 98.215 27.595 98.385 ;
        RECT 27.885 98.215 28.055 98.385 ;
        RECT 28.345 98.215 28.515 98.385 ;
        RECT 28.805 98.215 28.975 98.385 ;
        RECT 29.265 98.215 29.435 98.385 ;
        RECT 29.725 98.215 29.895 98.385 ;
        RECT 30.185 98.215 30.355 98.385 ;
        RECT 30.645 98.215 30.815 98.385 ;
        RECT 31.105 98.215 31.275 98.385 ;
        RECT 31.565 98.215 31.735 98.385 ;
        RECT 32.025 98.215 32.195 98.385 ;
        RECT 32.485 98.215 32.655 98.385 ;
        RECT 32.945 98.215 33.115 98.385 ;
        RECT 33.405 98.215 33.575 98.385 ;
        RECT 33.865 98.215 34.035 98.385 ;
        RECT 34.325 98.215 34.495 98.385 ;
        RECT 34.785 98.215 34.955 98.385 ;
        RECT 35.245 98.215 35.415 98.385 ;
        RECT 35.705 98.215 35.875 98.385 ;
        RECT 36.165 98.215 36.335 98.385 ;
        RECT 36.625 98.215 36.795 98.385 ;
        RECT 37.085 98.215 37.255 98.385 ;
        RECT 37.545 98.215 37.715 98.385 ;
        RECT 38.005 98.215 38.175 98.385 ;
        RECT 38.465 98.215 38.635 98.385 ;
        RECT 38.925 98.215 39.095 98.385 ;
        RECT 39.385 98.215 39.555 98.385 ;
        RECT 39.845 98.215 40.015 98.385 ;
        RECT 40.305 98.215 40.475 98.385 ;
        RECT 40.765 98.215 40.935 98.385 ;
        RECT 41.225 98.215 41.395 98.385 ;
        RECT 41.685 98.215 41.855 98.385 ;
        RECT 42.145 98.215 42.315 98.385 ;
        RECT 42.605 98.215 42.775 98.385 ;
        RECT 43.065 98.215 43.235 98.385 ;
        RECT 43.525 98.215 43.695 98.385 ;
        RECT 43.985 98.215 44.155 98.385 ;
        RECT 44.445 98.215 44.615 98.385 ;
        RECT 44.905 98.215 45.075 98.385 ;
        RECT 45.365 98.215 45.535 98.385 ;
        RECT 45.825 98.215 45.995 98.385 ;
        RECT 46.285 98.215 46.455 98.385 ;
        RECT 46.745 98.215 46.915 98.385 ;
        RECT 47.205 98.215 47.375 98.385 ;
        RECT 47.665 98.215 47.835 98.385 ;
        RECT 48.125 98.215 48.295 98.385 ;
        RECT 48.585 98.215 48.755 98.385 ;
        RECT 49.045 98.215 49.215 98.385 ;
        RECT 49.505 98.215 49.675 98.385 ;
        RECT 49.965 98.215 50.135 98.385 ;
        RECT 50.425 98.215 50.595 98.385 ;
        RECT 50.885 98.215 51.055 98.385 ;
        RECT 51.345 98.215 51.515 98.385 ;
        RECT 51.805 98.215 51.975 98.385 ;
        RECT 52.265 98.215 52.435 98.385 ;
        RECT 52.725 98.215 52.895 98.385 ;
        RECT 53.185 98.215 53.355 98.385 ;
        RECT 53.645 98.215 53.815 98.385 ;
        RECT 54.105 98.215 54.275 98.385 ;
        RECT 54.565 98.215 54.735 98.385 ;
        RECT 55.025 98.215 55.195 98.385 ;
        RECT 55.485 98.215 55.655 98.385 ;
        RECT 55.945 98.215 56.115 98.385 ;
        RECT 56.405 98.215 56.575 98.385 ;
        RECT 56.865 98.215 57.035 98.385 ;
        RECT 57.325 98.215 57.495 98.385 ;
        RECT 57.785 98.215 57.955 98.385 ;
        RECT 58.245 98.215 58.415 98.385 ;
        RECT 58.705 98.215 58.875 98.385 ;
        RECT 59.165 98.215 59.335 98.385 ;
        RECT 59.625 98.215 59.795 98.385 ;
        RECT 60.085 98.215 60.255 98.385 ;
        RECT 60.545 98.215 60.715 98.385 ;
        RECT 61.005 98.215 61.175 98.385 ;
        RECT 61.465 98.215 61.635 98.385 ;
        RECT 61.925 98.215 62.095 98.385 ;
        RECT 62.385 98.215 62.555 98.385 ;
        RECT 62.845 98.215 63.015 98.385 ;
        RECT 63.305 98.215 63.475 98.385 ;
        RECT 63.765 98.215 63.935 98.385 ;
        RECT 64.225 98.215 64.395 98.385 ;
        RECT 64.685 98.215 64.855 98.385 ;
        RECT 65.145 98.215 65.315 98.385 ;
        RECT 65.605 98.215 65.775 98.385 ;
        RECT 66.065 98.215 66.235 98.385 ;
        RECT 66.525 98.215 66.695 98.385 ;
        RECT 66.985 98.215 67.155 98.385 ;
        RECT 67.445 98.215 67.615 98.385 ;
        RECT 67.905 98.215 68.075 98.385 ;
        RECT 68.365 98.215 68.535 98.385 ;
        RECT 68.825 98.215 68.995 98.385 ;
        RECT 69.285 98.215 69.455 98.385 ;
        RECT 69.745 98.215 69.915 98.385 ;
        RECT 70.205 98.215 70.375 98.385 ;
        RECT 70.665 98.215 70.835 98.385 ;
        RECT 71.125 98.215 71.295 98.385 ;
        RECT 71.585 98.215 71.755 98.385 ;
        RECT 72.045 98.215 72.215 98.385 ;
        RECT 72.505 98.215 72.675 98.385 ;
        RECT 72.965 98.215 73.135 98.385 ;
        RECT 73.425 98.215 73.595 98.385 ;
        RECT 73.885 98.215 74.055 98.385 ;
        RECT 74.345 98.215 74.515 98.385 ;
        RECT 74.805 98.215 74.975 98.385 ;
        RECT 75.265 98.215 75.435 98.385 ;
        RECT 75.725 98.215 75.895 98.385 ;
        RECT 76.185 98.215 76.355 98.385 ;
        RECT 76.645 98.215 76.815 98.385 ;
        RECT 77.105 98.215 77.275 98.385 ;
        RECT 77.565 98.215 77.735 98.385 ;
        RECT 78.025 98.215 78.195 98.385 ;
        RECT 78.485 98.215 78.655 98.385 ;
        RECT 78.945 98.215 79.115 98.385 ;
        RECT 79.405 98.215 79.575 98.385 ;
        RECT 79.865 98.215 80.035 98.385 ;
        RECT 80.325 98.215 80.495 98.385 ;
        RECT 80.785 98.215 80.955 98.385 ;
        RECT 81.245 98.215 81.415 98.385 ;
        RECT 81.705 98.215 81.875 98.385 ;
        RECT 82.165 98.215 82.335 98.385 ;
        RECT 82.625 98.215 82.795 98.385 ;
        RECT 83.085 98.215 83.255 98.385 ;
        RECT 83.545 98.215 83.715 98.385 ;
        RECT 84.005 98.215 84.175 98.385 ;
        RECT 84.465 98.215 84.635 98.385 ;
        RECT 84.925 98.215 85.095 98.385 ;
        RECT 85.385 98.215 85.555 98.385 ;
        RECT 85.845 98.215 86.015 98.385 ;
        RECT 86.305 98.215 86.475 98.385 ;
        RECT 86.765 98.215 86.935 98.385 ;
        RECT 87.225 98.215 87.395 98.385 ;
        RECT 87.685 98.215 87.855 98.385 ;
        RECT 88.145 98.215 88.315 98.385 ;
        RECT 88.605 98.215 88.775 98.385 ;
        RECT 89.065 98.215 89.235 98.385 ;
        RECT 89.525 98.215 89.695 98.385 ;
        RECT 89.985 98.215 90.155 98.385 ;
        RECT 90.445 98.215 90.615 98.385 ;
        RECT 90.905 98.215 91.075 98.385 ;
        RECT 91.365 98.215 91.535 98.385 ;
        RECT 91.825 98.215 91.995 98.385 ;
        RECT 92.285 98.215 92.455 98.385 ;
        RECT 92.745 98.215 92.915 98.385 ;
        RECT 93.205 98.215 93.375 98.385 ;
        RECT 93.665 98.215 93.835 98.385 ;
        RECT 94.125 98.215 94.295 98.385 ;
        RECT 94.585 98.215 94.755 98.385 ;
        RECT 95.045 98.215 95.215 98.385 ;
        RECT 95.505 98.215 95.675 98.385 ;
        RECT 95.965 98.215 96.135 98.385 ;
        RECT 96.425 98.215 96.595 98.385 ;
        RECT 96.885 98.215 97.055 98.385 ;
        RECT 97.345 98.215 97.515 98.385 ;
        RECT 97.805 98.215 97.975 98.385 ;
        RECT 98.265 98.215 98.435 98.385 ;
        RECT 98.725 98.215 98.895 98.385 ;
        RECT 99.185 98.215 99.355 98.385 ;
        RECT 99.645 98.215 99.815 98.385 ;
        RECT 16.845 92.775 17.015 92.945 ;
        RECT 17.305 92.775 17.475 92.945 ;
        RECT 17.765 92.775 17.935 92.945 ;
        RECT 18.225 92.775 18.395 92.945 ;
        RECT 18.685 92.775 18.855 92.945 ;
        RECT 19.145 92.775 19.315 92.945 ;
        RECT 19.605 92.775 19.775 92.945 ;
        RECT 20.065 92.775 20.235 92.945 ;
        RECT 20.525 92.775 20.695 92.945 ;
        RECT 20.985 92.775 21.155 92.945 ;
        RECT 21.445 92.775 21.615 92.945 ;
        RECT 21.905 92.775 22.075 92.945 ;
        RECT 22.365 92.775 22.535 92.945 ;
        RECT 22.825 92.775 22.995 92.945 ;
        RECT 23.285 92.775 23.455 92.945 ;
        RECT 23.745 92.775 23.915 92.945 ;
        RECT 24.205 92.775 24.375 92.945 ;
        RECT 24.665 92.775 24.835 92.945 ;
        RECT 25.125 92.775 25.295 92.945 ;
        RECT 25.585 92.775 25.755 92.945 ;
        RECT 26.045 92.775 26.215 92.945 ;
        RECT 26.505 92.775 26.675 92.945 ;
        RECT 26.965 92.775 27.135 92.945 ;
        RECT 27.425 92.775 27.595 92.945 ;
        RECT 27.885 92.775 28.055 92.945 ;
        RECT 28.345 92.775 28.515 92.945 ;
        RECT 28.805 92.775 28.975 92.945 ;
        RECT 29.265 92.775 29.435 92.945 ;
        RECT 29.725 92.775 29.895 92.945 ;
        RECT 30.185 92.775 30.355 92.945 ;
        RECT 30.645 92.775 30.815 92.945 ;
        RECT 31.105 92.775 31.275 92.945 ;
        RECT 31.565 92.775 31.735 92.945 ;
        RECT 32.025 92.775 32.195 92.945 ;
        RECT 32.485 92.775 32.655 92.945 ;
        RECT 32.945 92.775 33.115 92.945 ;
        RECT 33.405 92.775 33.575 92.945 ;
        RECT 33.865 92.775 34.035 92.945 ;
        RECT 34.325 92.775 34.495 92.945 ;
        RECT 34.785 92.775 34.955 92.945 ;
        RECT 35.245 92.775 35.415 92.945 ;
        RECT 35.705 92.775 35.875 92.945 ;
        RECT 36.165 92.775 36.335 92.945 ;
        RECT 36.625 92.775 36.795 92.945 ;
        RECT 37.085 92.775 37.255 92.945 ;
        RECT 37.545 92.775 37.715 92.945 ;
        RECT 38.005 92.775 38.175 92.945 ;
        RECT 38.465 92.775 38.635 92.945 ;
        RECT 38.925 92.775 39.095 92.945 ;
        RECT 39.385 92.775 39.555 92.945 ;
        RECT 39.845 92.775 40.015 92.945 ;
        RECT 40.305 92.775 40.475 92.945 ;
        RECT 40.765 92.775 40.935 92.945 ;
        RECT 41.225 92.775 41.395 92.945 ;
        RECT 41.685 92.775 41.855 92.945 ;
        RECT 42.145 92.775 42.315 92.945 ;
        RECT 42.605 92.775 42.775 92.945 ;
        RECT 43.065 92.775 43.235 92.945 ;
        RECT 43.525 92.775 43.695 92.945 ;
        RECT 43.985 92.775 44.155 92.945 ;
        RECT 44.445 92.775 44.615 92.945 ;
        RECT 44.905 92.775 45.075 92.945 ;
        RECT 45.365 92.775 45.535 92.945 ;
        RECT 45.825 92.775 45.995 92.945 ;
        RECT 46.285 92.775 46.455 92.945 ;
        RECT 46.745 92.775 46.915 92.945 ;
        RECT 47.205 92.775 47.375 92.945 ;
        RECT 47.665 92.775 47.835 92.945 ;
        RECT 48.125 92.775 48.295 92.945 ;
        RECT 48.585 92.775 48.755 92.945 ;
        RECT 49.045 92.775 49.215 92.945 ;
        RECT 49.505 92.775 49.675 92.945 ;
        RECT 49.965 92.775 50.135 92.945 ;
        RECT 50.425 92.775 50.595 92.945 ;
        RECT 50.885 92.775 51.055 92.945 ;
        RECT 51.345 92.775 51.515 92.945 ;
        RECT 51.805 92.775 51.975 92.945 ;
        RECT 52.265 92.775 52.435 92.945 ;
        RECT 52.725 92.775 52.895 92.945 ;
        RECT 53.185 92.775 53.355 92.945 ;
        RECT 53.645 92.775 53.815 92.945 ;
        RECT 54.105 92.775 54.275 92.945 ;
        RECT 54.565 92.775 54.735 92.945 ;
        RECT 55.025 92.775 55.195 92.945 ;
        RECT 55.485 92.775 55.655 92.945 ;
        RECT 55.945 92.775 56.115 92.945 ;
        RECT 56.405 92.775 56.575 92.945 ;
        RECT 56.865 92.775 57.035 92.945 ;
        RECT 57.325 92.775 57.495 92.945 ;
        RECT 57.785 92.775 57.955 92.945 ;
        RECT 58.245 92.775 58.415 92.945 ;
        RECT 58.705 92.775 58.875 92.945 ;
        RECT 59.165 92.775 59.335 92.945 ;
        RECT 59.625 92.775 59.795 92.945 ;
        RECT 60.085 92.775 60.255 92.945 ;
        RECT 60.545 92.775 60.715 92.945 ;
        RECT 61.005 92.775 61.175 92.945 ;
        RECT 61.465 92.775 61.635 92.945 ;
        RECT 61.925 92.775 62.095 92.945 ;
        RECT 62.385 92.775 62.555 92.945 ;
        RECT 62.845 92.775 63.015 92.945 ;
        RECT 63.305 92.775 63.475 92.945 ;
        RECT 63.765 92.775 63.935 92.945 ;
        RECT 64.225 92.775 64.395 92.945 ;
        RECT 64.685 92.775 64.855 92.945 ;
        RECT 65.145 92.775 65.315 92.945 ;
        RECT 65.605 92.775 65.775 92.945 ;
        RECT 66.065 92.775 66.235 92.945 ;
        RECT 66.525 92.775 66.695 92.945 ;
        RECT 66.985 92.775 67.155 92.945 ;
        RECT 67.445 92.775 67.615 92.945 ;
        RECT 67.905 92.775 68.075 92.945 ;
        RECT 68.365 92.775 68.535 92.945 ;
        RECT 68.825 92.775 68.995 92.945 ;
        RECT 69.285 92.775 69.455 92.945 ;
        RECT 69.745 92.775 69.915 92.945 ;
        RECT 70.205 92.775 70.375 92.945 ;
        RECT 70.665 92.775 70.835 92.945 ;
        RECT 71.125 92.775 71.295 92.945 ;
        RECT 71.585 92.775 71.755 92.945 ;
        RECT 72.045 92.775 72.215 92.945 ;
        RECT 72.505 92.775 72.675 92.945 ;
        RECT 72.965 92.775 73.135 92.945 ;
        RECT 73.425 92.775 73.595 92.945 ;
        RECT 73.885 92.775 74.055 92.945 ;
        RECT 74.345 92.775 74.515 92.945 ;
        RECT 74.805 92.775 74.975 92.945 ;
        RECT 75.265 92.775 75.435 92.945 ;
        RECT 75.725 92.775 75.895 92.945 ;
        RECT 76.185 92.775 76.355 92.945 ;
        RECT 76.645 92.775 76.815 92.945 ;
        RECT 77.105 92.775 77.275 92.945 ;
        RECT 77.565 92.775 77.735 92.945 ;
        RECT 78.025 92.775 78.195 92.945 ;
        RECT 78.485 92.775 78.655 92.945 ;
        RECT 78.945 92.775 79.115 92.945 ;
        RECT 79.405 92.775 79.575 92.945 ;
        RECT 79.865 92.775 80.035 92.945 ;
        RECT 80.325 92.775 80.495 92.945 ;
        RECT 80.785 92.775 80.955 92.945 ;
        RECT 81.245 92.775 81.415 92.945 ;
        RECT 81.705 92.775 81.875 92.945 ;
        RECT 82.165 92.775 82.335 92.945 ;
        RECT 82.625 92.775 82.795 92.945 ;
        RECT 83.085 92.775 83.255 92.945 ;
        RECT 83.545 92.775 83.715 92.945 ;
        RECT 84.005 92.775 84.175 92.945 ;
        RECT 84.465 92.775 84.635 92.945 ;
        RECT 84.925 92.775 85.095 92.945 ;
        RECT 85.385 92.775 85.555 92.945 ;
        RECT 85.845 92.775 86.015 92.945 ;
        RECT 86.305 92.775 86.475 92.945 ;
        RECT 86.765 92.775 86.935 92.945 ;
        RECT 87.225 92.775 87.395 92.945 ;
        RECT 87.685 92.775 87.855 92.945 ;
        RECT 88.145 92.775 88.315 92.945 ;
        RECT 88.605 92.775 88.775 92.945 ;
        RECT 89.065 92.775 89.235 92.945 ;
        RECT 89.525 92.775 89.695 92.945 ;
        RECT 89.985 92.775 90.155 92.945 ;
        RECT 90.445 92.775 90.615 92.945 ;
        RECT 90.905 92.775 91.075 92.945 ;
        RECT 91.365 92.775 91.535 92.945 ;
        RECT 91.825 92.775 91.995 92.945 ;
        RECT 92.285 92.775 92.455 92.945 ;
        RECT 92.745 92.775 92.915 92.945 ;
        RECT 93.205 92.775 93.375 92.945 ;
        RECT 93.665 92.775 93.835 92.945 ;
        RECT 94.125 92.775 94.295 92.945 ;
        RECT 94.585 92.775 94.755 92.945 ;
        RECT 95.045 92.775 95.215 92.945 ;
        RECT 95.505 92.775 95.675 92.945 ;
        RECT 95.965 92.775 96.135 92.945 ;
        RECT 96.425 92.775 96.595 92.945 ;
        RECT 96.885 92.775 97.055 92.945 ;
        RECT 97.345 92.775 97.515 92.945 ;
        RECT 97.805 92.775 97.975 92.945 ;
        RECT 98.265 92.775 98.435 92.945 ;
        RECT 98.725 92.775 98.895 92.945 ;
        RECT 99.185 92.775 99.355 92.945 ;
        RECT 99.645 92.775 99.815 92.945 ;
        RECT 16.845 87.335 17.015 87.505 ;
        RECT 17.305 87.335 17.475 87.505 ;
        RECT 17.765 87.335 17.935 87.505 ;
        RECT 18.225 87.335 18.395 87.505 ;
        RECT 18.685 87.335 18.855 87.505 ;
        RECT 19.145 87.335 19.315 87.505 ;
        RECT 19.605 87.335 19.775 87.505 ;
        RECT 20.065 87.335 20.235 87.505 ;
        RECT 20.525 87.335 20.695 87.505 ;
        RECT 20.985 87.335 21.155 87.505 ;
        RECT 21.445 87.335 21.615 87.505 ;
        RECT 21.905 87.335 22.075 87.505 ;
        RECT 22.365 87.335 22.535 87.505 ;
        RECT 22.825 87.335 22.995 87.505 ;
        RECT 23.285 87.335 23.455 87.505 ;
        RECT 23.745 87.335 23.915 87.505 ;
        RECT 24.205 87.335 24.375 87.505 ;
        RECT 24.665 87.335 24.835 87.505 ;
        RECT 25.125 87.335 25.295 87.505 ;
        RECT 25.585 87.335 25.755 87.505 ;
        RECT 26.045 87.335 26.215 87.505 ;
        RECT 26.505 87.335 26.675 87.505 ;
        RECT 26.965 87.335 27.135 87.505 ;
        RECT 27.425 87.335 27.595 87.505 ;
        RECT 27.885 87.335 28.055 87.505 ;
        RECT 28.345 87.335 28.515 87.505 ;
        RECT 28.805 87.335 28.975 87.505 ;
        RECT 29.265 87.335 29.435 87.505 ;
        RECT 29.725 87.335 29.895 87.505 ;
        RECT 30.185 87.335 30.355 87.505 ;
        RECT 30.645 87.335 30.815 87.505 ;
        RECT 31.105 87.335 31.275 87.505 ;
        RECT 31.565 87.335 31.735 87.505 ;
        RECT 32.025 87.335 32.195 87.505 ;
        RECT 32.485 87.335 32.655 87.505 ;
        RECT 32.945 87.335 33.115 87.505 ;
        RECT 33.405 87.335 33.575 87.505 ;
        RECT 33.865 87.335 34.035 87.505 ;
        RECT 34.325 87.335 34.495 87.505 ;
        RECT 34.785 87.335 34.955 87.505 ;
        RECT 35.245 87.335 35.415 87.505 ;
        RECT 35.705 87.335 35.875 87.505 ;
        RECT 36.165 87.335 36.335 87.505 ;
        RECT 36.625 87.335 36.795 87.505 ;
        RECT 37.085 87.335 37.255 87.505 ;
        RECT 37.545 87.335 37.715 87.505 ;
        RECT 38.005 87.335 38.175 87.505 ;
        RECT 38.465 87.335 38.635 87.505 ;
        RECT 38.925 87.335 39.095 87.505 ;
        RECT 39.385 87.335 39.555 87.505 ;
        RECT 39.845 87.335 40.015 87.505 ;
        RECT 40.305 87.335 40.475 87.505 ;
        RECT 40.765 87.335 40.935 87.505 ;
        RECT 41.225 87.335 41.395 87.505 ;
        RECT 41.685 87.335 41.855 87.505 ;
        RECT 42.145 87.335 42.315 87.505 ;
        RECT 42.605 87.335 42.775 87.505 ;
        RECT 43.065 87.335 43.235 87.505 ;
        RECT 43.525 87.335 43.695 87.505 ;
        RECT 43.985 87.335 44.155 87.505 ;
        RECT 44.445 87.335 44.615 87.505 ;
        RECT 44.905 87.335 45.075 87.505 ;
        RECT 45.365 87.335 45.535 87.505 ;
        RECT 45.825 87.335 45.995 87.505 ;
        RECT 46.285 87.335 46.455 87.505 ;
        RECT 46.745 87.335 46.915 87.505 ;
        RECT 47.205 87.335 47.375 87.505 ;
        RECT 47.665 87.335 47.835 87.505 ;
        RECT 48.125 87.335 48.295 87.505 ;
        RECT 48.585 87.335 48.755 87.505 ;
        RECT 49.045 87.335 49.215 87.505 ;
        RECT 49.505 87.335 49.675 87.505 ;
        RECT 49.965 87.335 50.135 87.505 ;
        RECT 50.425 87.335 50.595 87.505 ;
        RECT 50.885 87.335 51.055 87.505 ;
        RECT 51.345 87.335 51.515 87.505 ;
        RECT 51.805 87.335 51.975 87.505 ;
        RECT 52.265 87.335 52.435 87.505 ;
        RECT 52.725 87.335 52.895 87.505 ;
        RECT 53.185 87.335 53.355 87.505 ;
        RECT 53.645 87.335 53.815 87.505 ;
        RECT 54.105 87.335 54.275 87.505 ;
        RECT 54.565 87.335 54.735 87.505 ;
        RECT 55.025 87.335 55.195 87.505 ;
        RECT 55.485 87.335 55.655 87.505 ;
        RECT 55.945 87.335 56.115 87.505 ;
        RECT 56.405 87.335 56.575 87.505 ;
        RECT 56.865 87.335 57.035 87.505 ;
        RECT 57.325 87.335 57.495 87.505 ;
        RECT 57.785 87.335 57.955 87.505 ;
        RECT 58.245 87.335 58.415 87.505 ;
        RECT 58.705 87.335 58.875 87.505 ;
        RECT 59.165 87.335 59.335 87.505 ;
        RECT 59.625 87.335 59.795 87.505 ;
        RECT 60.085 87.335 60.255 87.505 ;
        RECT 60.545 87.335 60.715 87.505 ;
        RECT 61.005 87.335 61.175 87.505 ;
        RECT 61.465 87.335 61.635 87.505 ;
        RECT 61.925 87.335 62.095 87.505 ;
        RECT 62.385 87.335 62.555 87.505 ;
        RECT 62.845 87.335 63.015 87.505 ;
        RECT 63.305 87.335 63.475 87.505 ;
        RECT 63.765 87.335 63.935 87.505 ;
        RECT 64.225 87.335 64.395 87.505 ;
        RECT 64.685 87.335 64.855 87.505 ;
        RECT 65.145 87.335 65.315 87.505 ;
        RECT 65.605 87.335 65.775 87.505 ;
        RECT 66.065 87.335 66.235 87.505 ;
        RECT 66.525 87.335 66.695 87.505 ;
        RECT 66.985 87.335 67.155 87.505 ;
        RECT 67.445 87.335 67.615 87.505 ;
        RECT 67.905 87.335 68.075 87.505 ;
        RECT 68.365 87.335 68.535 87.505 ;
        RECT 68.825 87.335 68.995 87.505 ;
        RECT 69.285 87.335 69.455 87.505 ;
        RECT 69.745 87.335 69.915 87.505 ;
        RECT 70.205 87.335 70.375 87.505 ;
        RECT 70.665 87.335 70.835 87.505 ;
        RECT 71.125 87.335 71.295 87.505 ;
        RECT 71.585 87.335 71.755 87.505 ;
        RECT 72.045 87.335 72.215 87.505 ;
        RECT 72.505 87.335 72.675 87.505 ;
        RECT 72.965 87.335 73.135 87.505 ;
        RECT 73.425 87.335 73.595 87.505 ;
        RECT 73.885 87.335 74.055 87.505 ;
        RECT 74.345 87.335 74.515 87.505 ;
        RECT 74.805 87.335 74.975 87.505 ;
        RECT 75.265 87.335 75.435 87.505 ;
        RECT 75.725 87.335 75.895 87.505 ;
        RECT 76.185 87.335 76.355 87.505 ;
        RECT 76.645 87.335 76.815 87.505 ;
        RECT 77.105 87.335 77.275 87.505 ;
        RECT 77.565 87.335 77.735 87.505 ;
        RECT 78.025 87.335 78.195 87.505 ;
        RECT 78.485 87.335 78.655 87.505 ;
        RECT 78.945 87.335 79.115 87.505 ;
        RECT 79.405 87.335 79.575 87.505 ;
        RECT 79.865 87.335 80.035 87.505 ;
        RECT 80.325 87.335 80.495 87.505 ;
        RECT 80.785 87.335 80.955 87.505 ;
        RECT 81.245 87.335 81.415 87.505 ;
        RECT 81.705 87.335 81.875 87.505 ;
        RECT 82.165 87.335 82.335 87.505 ;
        RECT 82.625 87.335 82.795 87.505 ;
        RECT 83.085 87.335 83.255 87.505 ;
        RECT 83.545 87.335 83.715 87.505 ;
        RECT 84.005 87.335 84.175 87.505 ;
        RECT 84.465 87.335 84.635 87.505 ;
        RECT 84.925 87.335 85.095 87.505 ;
        RECT 85.385 87.335 85.555 87.505 ;
        RECT 85.845 87.335 86.015 87.505 ;
        RECT 86.305 87.335 86.475 87.505 ;
        RECT 86.765 87.335 86.935 87.505 ;
        RECT 87.225 87.335 87.395 87.505 ;
        RECT 87.685 87.335 87.855 87.505 ;
        RECT 88.145 87.335 88.315 87.505 ;
        RECT 88.605 87.335 88.775 87.505 ;
        RECT 89.065 87.335 89.235 87.505 ;
        RECT 89.525 87.335 89.695 87.505 ;
        RECT 89.985 87.335 90.155 87.505 ;
        RECT 90.445 87.335 90.615 87.505 ;
        RECT 90.905 87.335 91.075 87.505 ;
        RECT 91.365 87.335 91.535 87.505 ;
        RECT 91.825 87.335 91.995 87.505 ;
        RECT 92.285 87.335 92.455 87.505 ;
        RECT 92.745 87.335 92.915 87.505 ;
        RECT 93.205 87.335 93.375 87.505 ;
        RECT 93.665 87.335 93.835 87.505 ;
        RECT 94.125 87.335 94.295 87.505 ;
        RECT 94.585 87.335 94.755 87.505 ;
        RECT 95.045 87.335 95.215 87.505 ;
        RECT 95.505 87.335 95.675 87.505 ;
        RECT 95.965 87.335 96.135 87.505 ;
        RECT 96.425 87.335 96.595 87.505 ;
        RECT 96.885 87.335 97.055 87.505 ;
        RECT 97.345 87.335 97.515 87.505 ;
        RECT 97.805 87.335 97.975 87.505 ;
        RECT 98.265 87.335 98.435 87.505 ;
        RECT 98.725 87.335 98.895 87.505 ;
        RECT 99.185 87.335 99.355 87.505 ;
        RECT 99.645 87.335 99.815 87.505 ;
        RECT 16.845 81.895 17.015 82.065 ;
        RECT 17.305 81.895 17.475 82.065 ;
        RECT 17.765 81.895 17.935 82.065 ;
        RECT 18.225 81.895 18.395 82.065 ;
        RECT 18.685 81.895 18.855 82.065 ;
        RECT 19.145 81.895 19.315 82.065 ;
        RECT 19.605 81.895 19.775 82.065 ;
        RECT 20.065 81.895 20.235 82.065 ;
        RECT 20.525 81.895 20.695 82.065 ;
        RECT 20.985 81.895 21.155 82.065 ;
        RECT 21.445 81.895 21.615 82.065 ;
        RECT 21.905 81.895 22.075 82.065 ;
        RECT 22.365 81.895 22.535 82.065 ;
        RECT 22.825 81.895 22.995 82.065 ;
        RECT 23.285 81.895 23.455 82.065 ;
        RECT 23.745 81.895 23.915 82.065 ;
        RECT 24.205 81.895 24.375 82.065 ;
        RECT 24.665 81.895 24.835 82.065 ;
        RECT 25.125 81.895 25.295 82.065 ;
        RECT 25.585 81.895 25.755 82.065 ;
        RECT 26.045 81.895 26.215 82.065 ;
        RECT 26.505 81.895 26.675 82.065 ;
        RECT 26.965 81.895 27.135 82.065 ;
        RECT 27.425 81.895 27.595 82.065 ;
        RECT 27.885 81.895 28.055 82.065 ;
        RECT 28.345 81.895 28.515 82.065 ;
        RECT 28.805 81.895 28.975 82.065 ;
        RECT 29.265 81.895 29.435 82.065 ;
        RECT 29.725 81.895 29.895 82.065 ;
        RECT 30.185 81.895 30.355 82.065 ;
        RECT 30.645 81.895 30.815 82.065 ;
        RECT 31.105 81.895 31.275 82.065 ;
        RECT 31.565 81.895 31.735 82.065 ;
        RECT 32.025 81.895 32.195 82.065 ;
        RECT 32.485 81.895 32.655 82.065 ;
        RECT 32.945 81.895 33.115 82.065 ;
        RECT 33.405 81.895 33.575 82.065 ;
        RECT 33.865 81.895 34.035 82.065 ;
        RECT 34.325 81.895 34.495 82.065 ;
        RECT 34.785 81.895 34.955 82.065 ;
        RECT 35.245 81.895 35.415 82.065 ;
        RECT 35.705 81.895 35.875 82.065 ;
        RECT 36.165 81.895 36.335 82.065 ;
        RECT 36.625 81.895 36.795 82.065 ;
        RECT 37.085 81.895 37.255 82.065 ;
        RECT 37.545 81.895 37.715 82.065 ;
        RECT 38.005 81.895 38.175 82.065 ;
        RECT 38.465 81.895 38.635 82.065 ;
        RECT 38.925 81.895 39.095 82.065 ;
        RECT 39.385 81.895 39.555 82.065 ;
        RECT 39.845 81.895 40.015 82.065 ;
        RECT 40.305 81.895 40.475 82.065 ;
        RECT 40.765 81.895 40.935 82.065 ;
        RECT 41.225 81.895 41.395 82.065 ;
        RECT 41.685 81.895 41.855 82.065 ;
        RECT 42.145 81.895 42.315 82.065 ;
        RECT 42.605 81.895 42.775 82.065 ;
        RECT 43.065 81.895 43.235 82.065 ;
        RECT 43.525 81.895 43.695 82.065 ;
        RECT 43.985 81.895 44.155 82.065 ;
        RECT 44.445 81.895 44.615 82.065 ;
        RECT 44.905 81.895 45.075 82.065 ;
        RECT 45.365 81.895 45.535 82.065 ;
        RECT 45.825 81.895 45.995 82.065 ;
        RECT 46.285 81.895 46.455 82.065 ;
        RECT 46.745 81.895 46.915 82.065 ;
        RECT 47.205 81.895 47.375 82.065 ;
        RECT 47.665 81.895 47.835 82.065 ;
        RECT 48.125 81.895 48.295 82.065 ;
        RECT 48.585 81.895 48.755 82.065 ;
        RECT 49.045 81.895 49.215 82.065 ;
        RECT 49.505 81.895 49.675 82.065 ;
        RECT 49.965 81.895 50.135 82.065 ;
        RECT 50.425 81.895 50.595 82.065 ;
        RECT 50.885 81.895 51.055 82.065 ;
        RECT 51.345 81.895 51.515 82.065 ;
        RECT 51.805 81.895 51.975 82.065 ;
        RECT 52.265 81.895 52.435 82.065 ;
        RECT 52.725 81.895 52.895 82.065 ;
        RECT 53.185 81.895 53.355 82.065 ;
        RECT 53.645 81.895 53.815 82.065 ;
        RECT 54.105 81.895 54.275 82.065 ;
        RECT 54.565 81.895 54.735 82.065 ;
        RECT 55.025 81.895 55.195 82.065 ;
        RECT 55.485 81.895 55.655 82.065 ;
        RECT 55.945 81.895 56.115 82.065 ;
        RECT 56.405 81.895 56.575 82.065 ;
        RECT 56.865 81.895 57.035 82.065 ;
        RECT 57.325 81.895 57.495 82.065 ;
        RECT 57.785 81.895 57.955 82.065 ;
        RECT 58.245 81.895 58.415 82.065 ;
        RECT 58.705 81.895 58.875 82.065 ;
        RECT 59.165 81.895 59.335 82.065 ;
        RECT 59.625 81.895 59.795 82.065 ;
        RECT 60.085 81.895 60.255 82.065 ;
        RECT 60.545 81.895 60.715 82.065 ;
        RECT 61.005 81.895 61.175 82.065 ;
        RECT 61.465 81.895 61.635 82.065 ;
        RECT 61.925 81.895 62.095 82.065 ;
        RECT 62.385 81.895 62.555 82.065 ;
        RECT 62.845 81.895 63.015 82.065 ;
        RECT 63.305 81.895 63.475 82.065 ;
        RECT 63.765 81.895 63.935 82.065 ;
        RECT 64.225 81.895 64.395 82.065 ;
        RECT 64.685 81.895 64.855 82.065 ;
        RECT 65.145 81.895 65.315 82.065 ;
        RECT 65.605 81.895 65.775 82.065 ;
        RECT 66.065 81.895 66.235 82.065 ;
        RECT 66.525 81.895 66.695 82.065 ;
        RECT 66.985 81.895 67.155 82.065 ;
        RECT 67.445 81.895 67.615 82.065 ;
        RECT 67.905 81.895 68.075 82.065 ;
        RECT 68.365 81.895 68.535 82.065 ;
        RECT 68.825 81.895 68.995 82.065 ;
        RECT 69.285 81.895 69.455 82.065 ;
        RECT 69.745 81.895 69.915 82.065 ;
        RECT 70.205 81.895 70.375 82.065 ;
        RECT 70.665 81.895 70.835 82.065 ;
        RECT 71.125 81.895 71.295 82.065 ;
        RECT 71.585 81.895 71.755 82.065 ;
        RECT 72.045 81.895 72.215 82.065 ;
        RECT 72.505 81.895 72.675 82.065 ;
        RECT 72.965 81.895 73.135 82.065 ;
        RECT 73.425 81.895 73.595 82.065 ;
        RECT 73.885 81.895 74.055 82.065 ;
        RECT 74.345 81.895 74.515 82.065 ;
        RECT 74.805 81.895 74.975 82.065 ;
        RECT 75.265 81.895 75.435 82.065 ;
        RECT 75.725 81.895 75.895 82.065 ;
        RECT 76.185 81.895 76.355 82.065 ;
        RECT 76.645 81.895 76.815 82.065 ;
        RECT 77.105 81.895 77.275 82.065 ;
        RECT 77.565 81.895 77.735 82.065 ;
        RECT 78.025 81.895 78.195 82.065 ;
        RECT 78.485 81.895 78.655 82.065 ;
        RECT 78.945 81.895 79.115 82.065 ;
        RECT 79.405 81.895 79.575 82.065 ;
        RECT 79.865 81.895 80.035 82.065 ;
        RECT 80.325 81.895 80.495 82.065 ;
        RECT 80.785 81.895 80.955 82.065 ;
        RECT 81.245 81.895 81.415 82.065 ;
        RECT 81.705 81.895 81.875 82.065 ;
        RECT 82.165 81.895 82.335 82.065 ;
        RECT 82.625 81.895 82.795 82.065 ;
        RECT 83.085 81.895 83.255 82.065 ;
        RECT 83.545 81.895 83.715 82.065 ;
        RECT 84.005 81.895 84.175 82.065 ;
        RECT 84.465 81.895 84.635 82.065 ;
        RECT 84.925 81.895 85.095 82.065 ;
        RECT 85.385 81.895 85.555 82.065 ;
        RECT 85.845 81.895 86.015 82.065 ;
        RECT 86.305 81.895 86.475 82.065 ;
        RECT 86.765 81.895 86.935 82.065 ;
        RECT 87.225 81.895 87.395 82.065 ;
        RECT 87.685 81.895 87.855 82.065 ;
        RECT 88.145 81.895 88.315 82.065 ;
        RECT 88.605 81.895 88.775 82.065 ;
        RECT 89.065 81.895 89.235 82.065 ;
        RECT 89.525 81.895 89.695 82.065 ;
        RECT 89.985 81.895 90.155 82.065 ;
        RECT 90.445 81.895 90.615 82.065 ;
        RECT 90.905 81.895 91.075 82.065 ;
        RECT 91.365 81.895 91.535 82.065 ;
        RECT 91.825 81.895 91.995 82.065 ;
        RECT 92.285 81.895 92.455 82.065 ;
        RECT 92.745 81.895 92.915 82.065 ;
        RECT 93.205 81.895 93.375 82.065 ;
        RECT 93.665 81.895 93.835 82.065 ;
        RECT 94.125 81.895 94.295 82.065 ;
        RECT 94.585 81.895 94.755 82.065 ;
        RECT 95.045 81.895 95.215 82.065 ;
        RECT 95.505 81.895 95.675 82.065 ;
        RECT 95.965 81.895 96.135 82.065 ;
        RECT 96.425 81.895 96.595 82.065 ;
        RECT 96.885 81.895 97.055 82.065 ;
        RECT 97.345 81.895 97.515 82.065 ;
        RECT 97.805 81.895 97.975 82.065 ;
        RECT 98.265 81.895 98.435 82.065 ;
        RECT 98.725 81.895 98.895 82.065 ;
        RECT 99.185 81.895 99.355 82.065 ;
        RECT 99.645 81.895 99.815 82.065 ;
        RECT 16.845 76.455 17.015 76.625 ;
        RECT 17.305 76.455 17.475 76.625 ;
        RECT 17.765 76.455 17.935 76.625 ;
        RECT 18.225 76.455 18.395 76.625 ;
        RECT 18.685 76.455 18.855 76.625 ;
        RECT 19.145 76.455 19.315 76.625 ;
        RECT 19.605 76.455 19.775 76.625 ;
        RECT 20.065 76.455 20.235 76.625 ;
        RECT 20.525 76.455 20.695 76.625 ;
        RECT 20.985 76.455 21.155 76.625 ;
        RECT 21.445 76.455 21.615 76.625 ;
        RECT 21.905 76.455 22.075 76.625 ;
        RECT 22.365 76.455 22.535 76.625 ;
        RECT 22.825 76.455 22.995 76.625 ;
        RECT 23.285 76.455 23.455 76.625 ;
        RECT 23.745 76.455 23.915 76.625 ;
        RECT 24.205 76.455 24.375 76.625 ;
        RECT 24.665 76.455 24.835 76.625 ;
        RECT 25.125 76.455 25.295 76.625 ;
        RECT 25.585 76.455 25.755 76.625 ;
        RECT 26.045 76.455 26.215 76.625 ;
        RECT 26.505 76.455 26.675 76.625 ;
        RECT 26.965 76.455 27.135 76.625 ;
        RECT 27.425 76.455 27.595 76.625 ;
        RECT 27.885 76.455 28.055 76.625 ;
        RECT 28.345 76.455 28.515 76.625 ;
        RECT 28.805 76.455 28.975 76.625 ;
        RECT 29.265 76.455 29.435 76.625 ;
        RECT 29.725 76.455 29.895 76.625 ;
        RECT 30.185 76.455 30.355 76.625 ;
        RECT 30.645 76.455 30.815 76.625 ;
        RECT 31.105 76.455 31.275 76.625 ;
        RECT 31.565 76.455 31.735 76.625 ;
        RECT 32.025 76.455 32.195 76.625 ;
        RECT 32.485 76.455 32.655 76.625 ;
        RECT 32.945 76.455 33.115 76.625 ;
        RECT 33.405 76.455 33.575 76.625 ;
        RECT 33.865 76.455 34.035 76.625 ;
        RECT 34.325 76.455 34.495 76.625 ;
        RECT 34.785 76.455 34.955 76.625 ;
        RECT 35.245 76.455 35.415 76.625 ;
        RECT 35.705 76.455 35.875 76.625 ;
        RECT 36.165 76.455 36.335 76.625 ;
        RECT 36.625 76.455 36.795 76.625 ;
        RECT 37.085 76.455 37.255 76.625 ;
        RECT 37.545 76.455 37.715 76.625 ;
        RECT 38.005 76.455 38.175 76.625 ;
        RECT 38.465 76.455 38.635 76.625 ;
        RECT 38.925 76.455 39.095 76.625 ;
        RECT 39.385 76.455 39.555 76.625 ;
        RECT 39.845 76.455 40.015 76.625 ;
        RECT 40.305 76.455 40.475 76.625 ;
        RECT 40.765 76.455 40.935 76.625 ;
        RECT 41.225 76.455 41.395 76.625 ;
        RECT 41.685 76.455 41.855 76.625 ;
        RECT 42.145 76.455 42.315 76.625 ;
        RECT 42.605 76.455 42.775 76.625 ;
        RECT 43.065 76.455 43.235 76.625 ;
        RECT 43.525 76.455 43.695 76.625 ;
        RECT 43.985 76.455 44.155 76.625 ;
        RECT 44.445 76.455 44.615 76.625 ;
        RECT 44.905 76.455 45.075 76.625 ;
        RECT 45.365 76.455 45.535 76.625 ;
        RECT 45.825 76.455 45.995 76.625 ;
        RECT 46.285 76.455 46.455 76.625 ;
        RECT 46.745 76.455 46.915 76.625 ;
        RECT 47.205 76.455 47.375 76.625 ;
        RECT 47.665 76.455 47.835 76.625 ;
        RECT 48.125 76.455 48.295 76.625 ;
        RECT 48.585 76.455 48.755 76.625 ;
        RECT 49.045 76.455 49.215 76.625 ;
        RECT 49.505 76.455 49.675 76.625 ;
        RECT 49.965 76.455 50.135 76.625 ;
        RECT 50.425 76.455 50.595 76.625 ;
        RECT 50.885 76.455 51.055 76.625 ;
        RECT 51.345 76.455 51.515 76.625 ;
        RECT 51.805 76.455 51.975 76.625 ;
        RECT 52.265 76.455 52.435 76.625 ;
        RECT 52.725 76.455 52.895 76.625 ;
        RECT 53.185 76.455 53.355 76.625 ;
        RECT 53.645 76.455 53.815 76.625 ;
        RECT 54.105 76.455 54.275 76.625 ;
        RECT 54.565 76.455 54.735 76.625 ;
        RECT 55.025 76.455 55.195 76.625 ;
        RECT 55.485 76.455 55.655 76.625 ;
        RECT 55.945 76.455 56.115 76.625 ;
        RECT 56.405 76.455 56.575 76.625 ;
        RECT 56.865 76.455 57.035 76.625 ;
        RECT 57.325 76.455 57.495 76.625 ;
        RECT 57.785 76.455 57.955 76.625 ;
        RECT 58.245 76.455 58.415 76.625 ;
        RECT 58.705 76.455 58.875 76.625 ;
        RECT 59.165 76.455 59.335 76.625 ;
        RECT 59.625 76.455 59.795 76.625 ;
        RECT 60.085 76.455 60.255 76.625 ;
        RECT 60.545 76.455 60.715 76.625 ;
        RECT 61.005 76.455 61.175 76.625 ;
        RECT 61.465 76.455 61.635 76.625 ;
        RECT 61.925 76.455 62.095 76.625 ;
        RECT 62.385 76.455 62.555 76.625 ;
        RECT 62.845 76.455 63.015 76.625 ;
        RECT 63.305 76.455 63.475 76.625 ;
        RECT 63.765 76.455 63.935 76.625 ;
        RECT 64.225 76.455 64.395 76.625 ;
        RECT 64.685 76.455 64.855 76.625 ;
        RECT 65.145 76.455 65.315 76.625 ;
        RECT 65.605 76.455 65.775 76.625 ;
        RECT 66.065 76.455 66.235 76.625 ;
        RECT 66.525 76.455 66.695 76.625 ;
        RECT 66.985 76.455 67.155 76.625 ;
        RECT 67.445 76.455 67.615 76.625 ;
        RECT 67.905 76.455 68.075 76.625 ;
        RECT 68.365 76.455 68.535 76.625 ;
        RECT 68.825 76.455 68.995 76.625 ;
        RECT 69.285 76.455 69.455 76.625 ;
        RECT 69.745 76.455 69.915 76.625 ;
        RECT 70.205 76.455 70.375 76.625 ;
        RECT 70.665 76.455 70.835 76.625 ;
        RECT 71.125 76.455 71.295 76.625 ;
        RECT 71.585 76.455 71.755 76.625 ;
        RECT 72.045 76.455 72.215 76.625 ;
        RECT 72.505 76.455 72.675 76.625 ;
        RECT 72.965 76.455 73.135 76.625 ;
        RECT 73.425 76.455 73.595 76.625 ;
        RECT 73.885 76.455 74.055 76.625 ;
        RECT 74.345 76.455 74.515 76.625 ;
        RECT 74.805 76.455 74.975 76.625 ;
        RECT 75.265 76.455 75.435 76.625 ;
        RECT 75.725 76.455 75.895 76.625 ;
        RECT 76.185 76.455 76.355 76.625 ;
        RECT 76.645 76.455 76.815 76.625 ;
        RECT 77.105 76.455 77.275 76.625 ;
        RECT 77.565 76.455 77.735 76.625 ;
        RECT 78.025 76.455 78.195 76.625 ;
        RECT 78.485 76.455 78.655 76.625 ;
        RECT 78.945 76.455 79.115 76.625 ;
        RECT 79.405 76.455 79.575 76.625 ;
        RECT 79.865 76.455 80.035 76.625 ;
        RECT 80.325 76.455 80.495 76.625 ;
        RECT 80.785 76.455 80.955 76.625 ;
        RECT 81.245 76.455 81.415 76.625 ;
        RECT 81.705 76.455 81.875 76.625 ;
        RECT 82.165 76.455 82.335 76.625 ;
        RECT 82.625 76.455 82.795 76.625 ;
        RECT 83.085 76.455 83.255 76.625 ;
        RECT 83.545 76.455 83.715 76.625 ;
        RECT 84.005 76.455 84.175 76.625 ;
        RECT 84.465 76.455 84.635 76.625 ;
        RECT 84.925 76.455 85.095 76.625 ;
        RECT 85.385 76.455 85.555 76.625 ;
        RECT 85.845 76.455 86.015 76.625 ;
        RECT 86.305 76.455 86.475 76.625 ;
        RECT 86.765 76.455 86.935 76.625 ;
        RECT 87.225 76.455 87.395 76.625 ;
        RECT 87.685 76.455 87.855 76.625 ;
        RECT 88.145 76.455 88.315 76.625 ;
        RECT 88.605 76.455 88.775 76.625 ;
        RECT 89.065 76.455 89.235 76.625 ;
        RECT 89.525 76.455 89.695 76.625 ;
        RECT 89.985 76.455 90.155 76.625 ;
        RECT 90.445 76.455 90.615 76.625 ;
        RECT 90.905 76.455 91.075 76.625 ;
        RECT 91.365 76.455 91.535 76.625 ;
        RECT 91.825 76.455 91.995 76.625 ;
        RECT 92.285 76.455 92.455 76.625 ;
        RECT 92.745 76.455 92.915 76.625 ;
        RECT 93.205 76.455 93.375 76.625 ;
        RECT 93.665 76.455 93.835 76.625 ;
        RECT 94.125 76.455 94.295 76.625 ;
        RECT 94.585 76.455 94.755 76.625 ;
        RECT 95.045 76.455 95.215 76.625 ;
        RECT 95.505 76.455 95.675 76.625 ;
        RECT 95.965 76.455 96.135 76.625 ;
        RECT 96.425 76.455 96.595 76.625 ;
        RECT 96.885 76.455 97.055 76.625 ;
        RECT 97.345 76.455 97.515 76.625 ;
        RECT 97.805 76.455 97.975 76.625 ;
        RECT 98.265 76.455 98.435 76.625 ;
        RECT 98.725 76.455 98.895 76.625 ;
        RECT 99.185 76.455 99.355 76.625 ;
        RECT 99.645 76.455 99.815 76.625 ;
        RECT 16.845 71.015 17.015 71.185 ;
        RECT 17.305 71.015 17.475 71.185 ;
        RECT 17.765 71.015 17.935 71.185 ;
        RECT 18.225 71.015 18.395 71.185 ;
        RECT 18.685 71.015 18.855 71.185 ;
        RECT 19.145 71.015 19.315 71.185 ;
        RECT 19.605 71.015 19.775 71.185 ;
        RECT 20.065 71.015 20.235 71.185 ;
        RECT 20.525 71.015 20.695 71.185 ;
        RECT 20.985 71.015 21.155 71.185 ;
        RECT 21.445 71.015 21.615 71.185 ;
        RECT 21.905 71.015 22.075 71.185 ;
        RECT 22.365 71.015 22.535 71.185 ;
        RECT 22.825 71.015 22.995 71.185 ;
        RECT 23.285 71.015 23.455 71.185 ;
        RECT 23.745 71.015 23.915 71.185 ;
        RECT 24.205 71.015 24.375 71.185 ;
        RECT 24.665 71.015 24.835 71.185 ;
        RECT 25.125 71.015 25.295 71.185 ;
        RECT 25.585 71.015 25.755 71.185 ;
        RECT 26.045 71.015 26.215 71.185 ;
        RECT 26.505 71.015 26.675 71.185 ;
        RECT 26.965 71.015 27.135 71.185 ;
        RECT 27.425 71.015 27.595 71.185 ;
        RECT 27.885 71.015 28.055 71.185 ;
        RECT 28.345 71.015 28.515 71.185 ;
        RECT 28.805 71.015 28.975 71.185 ;
        RECT 29.265 71.015 29.435 71.185 ;
        RECT 29.725 71.015 29.895 71.185 ;
        RECT 30.185 71.015 30.355 71.185 ;
        RECT 30.645 71.015 30.815 71.185 ;
        RECT 31.105 71.015 31.275 71.185 ;
        RECT 31.565 71.015 31.735 71.185 ;
        RECT 32.025 71.015 32.195 71.185 ;
        RECT 32.485 71.015 32.655 71.185 ;
        RECT 32.945 71.015 33.115 71.185 ;
        RECT 33.405 71.015 33.575 71.185 ;
        RECT 33.865 71.015 34.035 71.185 ;
        RECT 34.325 71.015 34.495 71.185 ;
        RECT 34.785 71.015 34.955 71.185 ;
        RECT 35.245 71.015 35.415 71.185 ;
        RECT 35.705 71.015 35.875 71.185 ;
        RECT 36.165 71.015 36.335 71.185 ;
        RECT 36.625 71.015 36.795 71.185 ;
        RECT 37.085 71.015 37.255 71.185 ;
        RECT 37.545 71.015 37.715 71.185 ;
        RECT 38.005 71.015 38.175 71.185 ;
        RECT 38.465 71.015 38.635 71.185 ;
        RECT 38.925 71.015 39.095 71.185 ;
        RECT 39.385 71.015 39.555 71.185 ;
        RECT 39.845 71.015 40.015 71.185 ;
        RECT 40.305 71.015 40.475 71.185 ;
        RECT 40.765 71.015 40.935 71.185 ;
        RECT 41.225 71.015 41.395 71.185 ;
        RECT 41.685 71.015 41.855 71.185 ;
        RECT 42.145 71.015 42.315 71.185 ;
        RECT 42.605 71.015 42.775 71.185 ;
        RECT 43.065 71.015 43.235 71.185 ;
        RECT 43.525 71.015 43.695 71.185 ;
        RECT 43.985 71.015 44.155 71.185 ;
        RECT 44.445 71.015 44.615 71.185 ;
        RECT 44.905 71.015 45.075 71.185 ;
        RECT 45.365 71.015 45.535 71.185 ;
        RECT 45.825 71.015 45.995 71.185 ;
        RECT 46.285 71.015 46.455 71.185 ;
        RECT 46.745 71.015 46.915 71.185 ;
        RECT 47.205 71.015 47.375 71.185 ;
        RECT 47.665 71.015 47.835 71.185 ;
        RECT 48.125 71.015 48.295 71.185 ;
        RECT 48.585 71.015 48.755 71.185 ;
        RECT 49.045 71.015 49.215 71.185 ;
        RECT 49.505 71.015 49.675 71.185 ;
        RECT 49.965 71.015 50.135 71.185 ;
        RECT 50.425 71.015 50.595 71.185 ;
        RECT 50.885 71.015 51.055 71.185 ;
        RECT 51.345 71.015 51.515 71.185 ;
        RECT 51.805 71.015 51.975 71.185 ;
        RECT 52.265 71.015 52.435 71.185 ;
        RECT 52.725 71.015 52.895 71.185 ;
        RECT 53.185 71.015 53.355 71.185 ;
        RECT 53.645 71.015 53.815 71.185 ;
        RECT 54.105 71.015 54.275 71.185 ;
        RECT 54.565 71.015 54.735 71.185 ;
        RECT 55.025 71.015 55.195 71.185 ;
        RECT 55.485 71.015 55.655 71.185 ;
        RECT 55.945 71.015 56.115 71.185 ;
        RECT 56.405 71.015 56.575 71.185 ;
        RECT 56.865 71.015 57.035 71.185 ;
        RECT 57.325 71.015 57.495 71.185 ;
        RECT 57.785 71.015 57.955 71.185 ;
        RECT 58.245 71.015 58.415 71.185 ;
        RECT 58.705 71.015 58.875 71.185 ;
        RECT 59.165 71.015 59.335 71.185 ;
        RECT 59.625 71.015 59.795 71.185 ;
        RECT 60.085 71.015 60.255 71.185 ;
        RECT 60.545 71.015 60.715 71.185 ;
        RECT 61.005 71.015 61.175 71.185 ;
        RECT 61.465 71.015 61.635 71.185 ;
        RECT 61.925 71.015 62.095 71.185 ;
        RECT 62.385 71.015 62.555 71.185 ;
        RECT 62.845 71.015 63.015 71.185 ;
        RECT 63.305 71.015 63.475 71.185 ;
        RECT 63.765 71.015 63.935 71.185 ;
        RECT 64.225 71.015 64.395 71.185 ;
        RECT 64.685 71.015 64.855 71.185 ;
        RECT 65.145 71.015 65.315 71.185 ;
        RECT 65.605 71.015 65.775 71.185 ;
        RECT 66.065 71.015 66.235 71.185 ;
        RECT 66.525 71.015 66.695 71.185 ;
        RECT 66.985 71.015 67.155 71.185 ;
        RECT 67.445 71.015 67.615 71.185 ;
        RECT 67.905 71.015 68.075 71.185 ;
        RECT 68.365 71.015 68.535 71.185 ;
        RECT 68.825 71.015 68.995 71.185 ;
        RECT 69.285 71.015 69.455 71.185 ;
        RECT 69.745 71.015 69.915 71.185 ;
        RECT 70.205 71.015 70.375 71.185 ;
        RECT 70.665 71.015 70.835 71.185 ;
        RECT 71.125 71.015 71.295 71.185 ;
        RECT 71.585 71.015 71.755 71.185 ;
        RECT 72.045 71.015 72.215 71.185 ;
        RECT 72.505 71.015 72.675 71.185 ;
        RECT 72.965 71.015 73.135 71.185 ;
        RECT 73.425 71.015 73.595 71.185 ;
        RECT 73.885 71.015 74.055 71.185 ;
        RECT 74.345 71.015 74.515 71.185 ;
        RECT 74.805 71.015 74.975 71.185 ;
        RECT 75.265 71.015 75.435 71.185 ;
        RECT 75.725 71.015 75.895 71.185 ;
        RECT 76.185 71.015 76.355 71.185 ;
        RECT 76.645 71.015 76.815 71.185 ;
        RECT 77.105 71.015 77.275 71.185 ;
        RECT 77.565 71.015 77.735 71.185 ;
        RECT 78.025 71.015 78.195 71.185 ;
        RECT 78.485 71.015 78.655 71.185 ;
        RECT 78.945 71.015 79.115 71.185 ;
        RECT 79.405 71.015 79.575 71.185 ;
        RECT 79.865 71.015 80.035 71.185 ;
        RECT 80.325 71.015 80.495 71.185 ;
        RECT 80.785 71.015 80.955 71.185 ;
        RECT 81.245 71.015 81.415 71.185 ;
        RECT 81.705 71.015 81.875 71.185 ;
        RECT 82.165 71.015 82.335 71.185 ;
        RECT 82.625 71.015 82.795 71.185 ;
        RECT 83.085 71.015 83.255 71.185 ;
        RECT 83.545 71.015 83.715 71.185 ;
        RECT 84.005 71.015 84.175 71.185 ;
        RECT 84.465 71.015 84.635 71.185 ;
        RECT 84.925 71.015 85.095 71.185 ;
        RECT 85.385 71.015 85.555 71.185 ;
        RECT 85.845 71.015 86.015 71.185 ;
        RECT 86.305 71.015 86.475 71.185 ;
        RECT 86.765 71.015 86.935 71.185 ;
        RECT 87.225 71.015 87.395 71.185 ;
        RECT 87.685 71.015 87.855 71.185 ;
        RECT 88.145 71.015 88.315 71.185 ;
        RECT 88.605 71.015 88.775 71.185 ;
        RECT 89.065 71.015 89.235 71.185 ;
        RECT 89.525 71.015 89.695 71.185 ;
        RECT 89.985 71.015 90.155 71.185 ;
        RECT 90.445 71.015 90.615 71.185 ;
        RECT 90.905 71.015 91.075 71.185 ;
        RECT 91.365 71.015 91.535 71.185 ;
        RECT 91.825 71.015 91.995 71.185 ;
        RECT 92.285 71.015 92.455 71.185 ;
        RECT 92.745 71.015 92.915 71.185 ;
        RECT 93.205 71.015 93.375 71.185 ;
        RECT 93.665 71.015 93.835 71.185 ;
        RECT 94.125 71.015 94.295 71.185 ;
        RECT 94.585 71.015 94.755 71.185 ;
        RECT 95.045 71.015 95.215 71.185 ;
        RECT 95.505 71.015 95.675 71.185 ;
        RECT 95.965 71.015 96.135 71.185 ;
        RECT 96.425 71.015 96.595 71.185 ;
        RECT 96.885 71.015 97.055 71.185 ;
        RECT 97.345 71.015 97.515 71.185 ;
        RECT 97.805 71.015 97.975 71.185 ;
        RECT 98.265 71.015 98.435 71.185 ;
        RECT 98.725 71.015 98.895 71.185 ;
        RECT 99.185 71.015 99.355 71.185 ;
        RECT 99.645 71.015 99.815 71.185 ;
        RECT 16.845 65.575 17.015 65.745 ;
        RECT 17.305 65.575 17.475 65.745 ;
        RECT 17.765 65.575 17.935 65.745 ;
        RECT 18.225 65.575 18.395 65.745 ;
        RECT 18.685 65.575 18.855 65.745 ;
        RECT 19.145 65.575 19.315 65.745 ;
        RECT 19.605 65.575 19.775 65.745 ;
        RECT 20.065 65.575 20.235 65.745 ;
        RECT 20.525 65.575 20.695 65.745 ;
        RECT 20.985 65.575 21.155 65.745 ;
        RECT 21.445 65.575 21.615 65.745 ;
        RECT 21.905 65.575 22.075 65.745 ;
        RECT 22.365 65.575 22.535 65.745 ;
        RECT 22.825 65.575 22.995 65.745 ;
        RECT 23.285 65.575 23.455 65.745 ;
        RECT 23.745 65.575 23.915 65.745 ;
        RECT 24.205 65.575 24.375 65.745 ;
        RECT 24.665 65.575 24.835 65.745 ;
        RECT 25.125 65.575 25.295 65.745 ;
        RECT 25.585 65.575 25.755 65.745 ;
        RECT 26.045 65.575 26.215 65.745 ;
        RECT 26.505 65.575 26.675 65.745 ;
        RECT 26.965 65.575 27.135 65.745 ;
        RECT 27.425 65.575 27.595 65.745 ;
        RECT 27.885 65.575 28.055 65.745 ;
        RECT 28.345 65.575 28.515 65.745 ;
        RECT 28.805 65.575 28.975 65.745 ;
        RECT 29.265 65.575 29.435 65.745 ;
        RECT 29.725 65.575 29.895 65.745 ;
        RECT 30.185 65.575 30.355 65.745 ;
        RECT 30.645 65.575 30.815 65.745 ;
        RECT 31.105 65.575 31.275 65.745 ;
        RECT 31.565 65.575 31.735 65.745 ;
        RECT 32.025 65.575 32.195 65.745 ;
        RECT 32.485 65.575 32.655 65.745 ;
        RECT 32.945 65.575 33.115 65.745 ;
        RECT 33.405 65.575 33.575 65.745 ;
        RECT 33.865 65.575 34.035 65.745 ;
        RECT 34.325 65.575 34.495 65.745 ;
        RECT 34.785 65.575 34.955 65.745 ;
        RECT 35.245 65.575 35.415 65.745 ;
        RECT 35.705 65.575 35.875 65.745 ;
        RECT 36.165 65.575 36.335 65.745 ;
        RECT 36.625 65.575 36.795 65.745 ;
        RECT 37.085 65.575 37.255 65.745 ;
        RECT 37.545 65.575 37.715 65.745 ;
        RECT 38.005 65.575 38.175 65.745 ;
        RECT 38.465 65.575 38.635 65.745 ;
        RECT 38.925 65.575 39.095 65.745 ;
        RECT 39.385 65.575 39.555 65.745 ;
        RECT 39.845 65.575 40.015 65.745 ;
        RECT 40.305 65.575 40.475 65.745 ;
        RECT 40.765 65.575 40.935 65.745 ;
        RECT 41.225 65.575 41.395 65.745 ;
        RECT 41.685 65.575 41.855 65.745 ;
        RECT 42.145 65.575 42.315 65.745 ;
        RECT 42.605 65.575 42.775 65.745 ;
        RECT 43.065 65.575 43.235 65.745 ;
        RECT 43.525 65.575 43.695 65.745 ;
        RECT 43.985 65.575 44.155 65.745 ;
        RECT 44.445 65.575 44.615 65.745 ;
        RECT 44.905 65.575 45.075 65.745 ;
        RECT 45.365 65.575 45.535 65.745 ;
        RECT 45.825 65.575 45.995 65.745 ;
        RECT 46.285 65.575 46.455 65.745 ;
        RECT 46.745 65.575 46.915 65.745 ;
        RECT 47.205 65.575 47.375 65.745 ;
        RECT 47.665 65.575 47.835 65.745 ;
        RECT 48.125 65.575 48.295 65.745 ;
        RECT 48.585 65.575 48.755 65.745 ;
        RECT 49.045 65.575 49.215 65.745 ;
        RECT 49.505 65.575 49.675 65.745 ;
        RECT 49.965 65.575 50.135 65.745 ;
        RECT 50.425 65.575 50.595 65.745 ;
        RECT 50.885 65.575 51.055 65.745 ;
        RECT 51.345 65.575 51.515 65.745 ;
        RECT 51.805 65.575 51.975 65.745 ;
        RECT 52.265 65.575 52.435 65.745 ;
        RECT 52.725 65.575 52.895 65.745 ;
        RECT 53.185 65.575 53.355 65.745 ;
        RECT 53.645 65.575 53.815 65.745 ;
        RECT 54.105 65.575 54.275 65.745 ;
        RECT 54.565 65.575 54.735 65.745 ;
        RECT 55.025 65.575 55.195 65.745 ;
        RECT 55.485 65.575 55.655 65.745 ;
        RECT 55.945 65.575 56.115 65.745 ;
        RECT 56.405 65.575 56.575 65.745 ;
        RECT 56.865 65.575 57.035 65.745 ;
        RECT 57.325 65.575 57.495 65.745 ;
        RECT 57.785 65.575 57.955 65.745 ;
        RECT 58.245 65.575 58.415 65.745 ;
        RECT 58.705 65.575 58.875 65.745 ;
        RECT 59.165 65.575 59.335 65.745 ;
        RECT 59.625 65.575 59.795 65.745 ;
        RECT 60.085 65.575 60.255 65.745 ;
        RECT 60.545 65.575 60.715 65.745 ;
        RECT 61.005 65.575 61.175 65.745 ;
        RECT 61.465 65.575 61.635 65.745 ;
        RECT 61.925 65.575 62.095 65.745 ;
        RECT 62.385 65.575 62.555 65.745 ;
        RECT 62.845 65.575 63.015 65.745 ;
        RECT 63.305 65.575 63.475 65.745 ;
        RECT 63.765 65.575 63.935 65.745 ;
        RECT 64.225 65.575 64.395 65.745 ;
        RECT 64.685 65.575 64.855 65.745 ;
        RECT 65.145 65.575 65.315 65.745 ;
        RECT 65.605 65.575 65.775 65.745 ;
        RECT 66.065 65.575 66.235 65.745 ;
        RECT 66.525 65.575 66.695 65.745 ;
        RECT 66.985 65.575 67.155 65.745 ;
        RECT 67.445 65.575 67.615 65.745 ;
        RECT 67.905 65.575 68.075 65.745 ;
        RECT 68.365 65.575 68.535 65.745 ;
        RECT 68.825 65.575 68.995 65.745 ;
        RECT 69.285 65.575 69.455 65.745 ;
        RECT 69.745 65.575 69.915 65.745 ;
        RECT 70.205 65.575 70.375 65.745 ;
        RECT 70.665 65.575 70.835 65.745 ;
        RECT 71.125 65.575 71.295 65.745 ;
        RECT 71.585 65.575 71.755 65.745 ;
        RECT 72.045 65.575 72.215 65.745 ;
        RECT 72.505 65.575 72.675 65.745 ;
        RECT 72.965 65.575 73.135 65.745 ;
        RECT 73.425 65.575 73.595 65.745 ;
        RECT 73.885 65.575 74.055 65.745 ;
        RECT 74.345 65.575 74.515 65.745 ;
        RECT 74.805 65.575 74.975 65.745 ;
        RECT 75.265 65.575 75.435 65.745 ;
        RECT 75.725 65.575 75.895 65.745 ;
        RECT 76.185 65.575 76.355 65.745 ;
        RECT 76.645 65.575 76.815 65.745 ;
        RECT 77.105 65.575 77.275 65.745 ;
        RECT 77.565 65.575 77.735 65.745 ;
        RECT 78.025 65.575 78.195 65.745 ;
        RECT 78.485 65.575 78.655 65.745 ;
        RECT 78.945 65.575 79.115 65.745 ;
        RECT 79.405 65.575 79.575 65.745 ;
        RECT 79.865 65.575 80.035 65.745 ;
        RECT 80.325 65.575 80.495 65.745 ;
        RECT 80.785 65.575 80.955 65.745 ;
        RECT 81.245 65.575 81.415 65.745 ;
        RECT 81.705 65.575 81.875 65.745 ;
        RECT 82.165 65.575 82.335 65.745 ;
        RECT 82.625 65.575 82.795 65.745 ;
        RECT 83.085 65.575 83.255 65.745 ;
        RECT 83.545 65.575 83.715 65.745 ;
        RECT 84.005 65.575 84.175 65.745 ;
        RECT 84.465 65.575 84.635 65.745 ;
        RECT 84.925 65.575 85.095 65.745 ;
        RECT 85.385 65.575 85.555 65.745 ;
        RECT 85.845 65.575 86.015 65.745 ;
        RECT 86.305 65.575 86.475 65.745 ;
        RECT 86.765 65.575 86.935 65.745 ;
        RECT 87.225 65.575 87.395 65.745 ;
        RECT 87.685 65.575 87.855 65.745 ;
        RECT 88.145 65.575 88.315 65.745 ;
        RECT 88.605 65.575 88.775 65.745 ;
        RECT 89.065 65.575 89.235 65.745 ;
        RECT 89.525 65.575 89.695 65.745 ;
        RECT 89.985 65.575 90.155 65.745 ;
        RECT 90.445 65.575 90.615 65.745 ;
        RECT 90.905 65.575 91.075 65.745 ;
        RECT 91.365 65.575 91.535 65.745 ;
        RECT 91.825 65.575 91.995 65.745 ;
        RECT 92.285 65.575 92.455 65.745 ;
        RECT 92.745 65.575 92.915 65.745 ;
        RECT 93.205 65.575 93.375 65.745 ;
        RECT 93.665 65.575 93.835 65.745 ;
        RECT 94.125 65.575 94.295 65.745 ;
        RECT 94.585 65.575 94.755 65.745 ;
        RECT 95.045 65.575 95.215 65.745 ;
        RECT 95.505 65.575 95.675 65.745 ;
        RECT 95.965 65.575 96.135 65.745 ;
        RECT 96.425 65.575 96.595 65.745 ;
        RECT 96.885 65.575 97.055 65.745 ;
        RECT 97.345 65.575 97.515 65.745 ;
        RECT 97.805 65.575 97.975 65.745 ;
        RECT 98.265 65.575 98.435 65.745 ;
        RECT 98.725 65.575 98.895 65.745 ;
        RECT 99.185 65.575 99.355 65.745 ;
        RECT 99.645 65.575 99.815 65.745 ;
        RECT 16.845 60.135 17.015 60.305 ;
        RECT 17.305 60.135 17.475 60.305 ;
        RECT 17.765 60.135 17.935 60.305 ;
        RECT 18.225 60.135 18.395 60.305 ;
        RECT 18.685 60.135 18.855 60.305 ;
        RECT 19.145 60.135 19.315 60.305 ;
        RECT 19.605 60.135 19.775 60.305 ;
        RECT 20.065 60.135 20.235 60.305 ;
        RECT 20.525 60.135 20.695 60.305 ;
        RECT 20.985 60.135 21.155 60.305 ;
        RECT 21.445 60.135 21.615 60.305 ;
        RECT 21.905 60.135 22.075 60.305 ;
        RECT 22.365 60.135 22.535 60.305 ;
        RECT 22.825 60.135 22.995 60.305 ;
        RECT 23.285 60.135 23.455 60.305 ;
        RECT 23.745 60.135 23.915 60.305 ;
        RECT 24.205 60.135 24.375 60.305 ;
        RECT 24.665 60.135 24.835 60.305 ;
        RECT 25.125 60.135 25.295 60.305 ;
        RECT 25.585 60.135 25.755 60.305 ;
        RECT 26.045 60.135 26.215 60.305 ;
        RECT 26.505 60.135 26.675 60.305 ;
        RECT 26.965 60.135 27.135 60.305 ;
        RECT 27.425 60.135 27.595 60.305 ;
        RECT 27.885 60.135 28.055 60.305 ;
        RECT 28.345 60.135 28.515 60.305 ;
        RECT 28.805 60.135 28.975 60.305 ;
        RECT 29.265 60.135 29.435 60.305 ;
        RECT 29.725 60.135 29.895 60.305 ;
        RECT 30.185 60.135 30.355 60.305 ;
        RECT 30.645 60.135 30.815 60.305 ;
        RECT 31.105 60.135 31.275 60.305 ;
        RECT 31.565 60.135 31.735 60.305 ;
        RECT 32.025 60.135 32.195 60.305 ;
        RECT 32.485 60.135 32.655 60.305 ;
        RECT 32.945 60.135 33.115 60.305 ;
        RECT 33.405 60.135 33.575 60.305 ;
        RECT 33.865 60.135 34.035 60.305 ;
        RECT 34.325 60.135 34.495 60.305 ;
        RECT 34.785 60.135 34.955 60.305 ;
        RECT 35.245 60.135 35.415 60.305 ;
        RECT 35.705 60.135 35.875 60.305 ;
        RECT 36.165 60.135 36.335 60.305 ;
        RECT 36.625 60.135 36.795 60.305 ;
        RECT 37.085 60.135 37.255 60.305 ;
        RECT 37.545 60.135 37.715 60.305 ;
        RECT 38.005 60.135 38.175 60.305 ;
        RECT 38.465 60.135 38.635 60.305 ;
        RECT 38.925 60.135 39.095 60.305 ;
        RECT 39.385 60.135 39.555 60.305 ;
        RECT 39.845 60.135 40.015 60.305 ;
        RECT 40.305 60.135 40.475 60.305 ;
        RECT 40.765 60.135 40.935 60.305 ;
        RECT 41.225 60.135 41.395 60.305 ;
        RECT 41.685 60.135 41.855 60.305 ;
        RECT 42.145 60.135 42.315 60.305 ;
        RECT 42.605 60.135 42.775 60.305 ;
        RECT 43.065 60.135 43.235 60.305 ;
        RECT 43.525 60.135 43.695 60.305 ;
        RECT 43.985 60.135 44.155 60.305 ;
        RECT 44.445 60.135 44.615 60.305 ;
        RECT 44.905 60.135 45.075 60.305 ;
        RECT 45.365 60.135 45.535 60.305 ;
        RECT 45.825 60.135 45.995 60.305 ;
        RECT 46.285 60.135 46.455 60.305 ;
        RECT 46.745 60.135 46.915 60.305 ;
        RECT 47.205 60.135 47.375 60.305 ;
        RECT 47.665 60.135 47.835 60.305 ;
        RECT 48.125 60.135 48.295 60.305 ;
        RECT 48.585 60.135 48.755 60.305 ;
        RECT 49.045 60.135 49.215 60.305 ;
        RECT 49.505 60.135 49.675 60.305 ;
        RECT 49.965 60.135 50.135 60.305 ;
        RECT 50.425 60.135 50.595 60.305 ;
        RECT 50.885 60.135 51.055 60.305 ;
        RECT 51.345 60.135 51.515 60.305 ;
        RECT 51.805 60.135 51.975 60.305 ;
        RECT 52.265 60.135 52.435 60.305 ;
        RECT 52.725 60.135 52.895 60.305 ;
        RECT 53.185 60.135 53.355 60.305 ;
        RECT 53.645 60.135 53.815 60.305 ;
        RECT 54.105 60.135 54.275 60.305 ;
        RECT 54.565 60.135 54.735 60.305 ;
        RECT 55.025 60.135 55.195 60.305 ;
        RECT 55.485 60.135 55.655 60.305 ;
        RECT 55.945 60.135 56.115 60.305 ;
        RECT 56.405 60.135 56.575 60.305 ;
        RECT 56.865 60.135 57.035 60.305 ;
        RECT 57.325 60.135 57.495 60.305 ;
        RECT 57.785 60.135 57.955 60.305 ;
        RECT 58.245 60.135 58.415 60.305 ;
        RECT 58.705 60.135 58.875 60.305 ;
        RECT 59.165 60.135 59.335 60.305 ;
        RECT 59.625 60.135 59.795 60.305 ;
        RECT 60.085 60.135 60.255 60.305 ;
        RECT 60.545 60.135 60.715 60.305 ;
        RECT 61.005 60.135 61.175 60.305 ;
        RECT 61.465 60.135 61.635 60.305 ;
        RECT 61.925 60.135 62.095 60.305 ;
        RECT 62.385 60.135 62.555 60.305 ;
        RECT 62.845 60.135 63.015 60.305 ;
        RECT 63.305 60.135 63.475 60.305 ;
        RECT 63.765 60.135 63.935 60.305 ;
        RECT 64.225 60.135 64.395 60.305 ;
        RECT 64.685 60.135 64.855 60.305 ;
        RECT 65.145 60.135 65.315 60.305 ;
        RECT 65.605 60.135 65.775 60.305 ;
        RECT 66.065 60.135 66.235 60.305 ;
        RECT 66.525 60.135 66.695 60.305 ;
        RECT 66.985 60.135 67.155 60.305 ;
        RECT 67.445 60.135 67.615 60.305 ;
        RECT 67.905 60.135 68.075 60.305 ;
        RECT 68.365 60.135 68.535 60.305 ;
        RECT 68.825 60.135 68.995 60.305 ;
        RECT 69.285 60.135 69.455 60.305 ;
        RECT 69.745 60.135 69.915 60.305 ;
        RECT 70.205 60.135 70.375 60.305 ;
        RECT 70.665 60.135 70.835 60.305 ;
        RECT 71.125 60.135 71.295 60.305 ;
        RECT 71.585 60.135 71.755 60.305 ;
        RECT 72.045 60.135 72.215 60.305 ;
        RECT 72.505 60.135 72.675 60.305 ;
        RECT 72.965 60.135 73.135 60.305 ;
        RECT 73.425 60.135 73.595 60.305 ;
        RECT 73.885 60.135 74.055 60.305 ;
        RECT 74.345 60.135 74.515 60.305 ;
        RECT 74.805 60.135 74.975 60.305 ;
        RECT 75.265 60.135 75.435 60.305 ;
        RECT 75.725 60.135 75.895 60.305 ;
        RECT 76.185 60.135 76.355 60.305 ;
        RECT 76.645 60.135 76.815 60.305 ;
        RECT 77.105 60.135 77.275 60.305 ;
        RECT 77.565 60.135 77.735 60.305 ;
        RECT 78.025 60.135 78.195 60.305 ;
        RECT 78.485 60.135 78.655 60.305 ;
        RECT 78.945 60.135 79.115 60.305 ;
        RECT 79.405 60.135 79.575 60.305 ;
        RECT 79.865 60.135 80.035 60.305 ;
        RECT 80.325 60.135 80.495 60.305 ;
        RECT 80.785 60.135 80.955 60.305 ;
        RECT 81.245 60.135 81.415 60.305 ;
        RECT 81.705 60.135 81.875 60.305 ;
        RECT 82.165 60.135 82.335 60.305 ;
        RECT 82.625 60.135 82.795 60.305 ;
        RECT 83.085 60.135 83.255 60.305 ;
        RECT 83.545 60.135 83.715 60.305 ;
        RECT 84.005 60.135 84.175 60.305 ;
        RECT 84.465 60.135 84.635 60.305 ;
        RECT 84.925 60.135 85.095 60.305 ;
        RECT 85.385 60.135 85.555 60.305 ;
        RECT 85.845 60.135 86.015 60.305 ;
        RECT 86.305 60.135 86.475 60.305 ;
        RECT 86.765 60.135 86.935 60.305 ;
        RECT 87.225 60.135 87.395 60.305 ;
        RECT 87.685 60.135 87.855 60.305 ;
        RECT 88.145 60.135 88.315 60.305 ;
        RECT 88.605 60.135 88.775 60.305 ;
        RECT 89.065 60.135 89.235 60.305 ;
        RECT 89.525 60.135 89.695 60.305 ;
        RECT 89.985 60.135 90.155 60.305 ;
        RECT 90.445 60.135 90.615 60.305 ;
        RECT 90.905 60.135 91.075 60.305 ;
        RECT 91.365 60.135 91.535 60.305 ;
        RECT 91.825 60.135 91.995 60.305 ;
        RECT 92.285 60.135 92.455 60.305 ;
        RECT 92.745 60.135 92.915 60.305 ;
        RECT 93.205 60.135 93.375 60.305 ;
        RECT 93.665 60.135 93.835 60.305 ;
        RECT 94.125 60.135 94.295 60.305 ;
        RECT 94.585 60.135 94.755 60.305 ;
        RECT 95.045 60.135 95.215 60.305 ;
        RECT 95.505 60.135 95.675 60.305 ;
        RECT 95.965 60.135 96.135 60.305 ;
        RECT 96.425 60.135 96.595 60.305 ;
        RECT 96.885 60.135 97.055 60.305 ;
        RECT 97.345 60.135 97.515 60.305 ;
        RECT 97.805 60.135 97.975 60.305 ;
        RECT 98.265 60.135 98.435 60.305 ;
        RECT 98.725 60.135 98.895 60.305 ;
        RECT 99.185 60.135 99.355 60.305 ;
        RECT 99.645 60.135 99.815 60.305 ;
        RECT 16.845 54.695 17.015 54.865 ;
        RECT 17.305 54.695 17.475 54.865 ;
        RECT 17.765 54.695 17.935 54.865 ;
        RECT 18.225 54.695 18.395 54.865 ;
        RECT 18.685 54.695 18.855 54.865 ;
        RECT 19.145 54.695 19.315 54.865 ;
        RECT 19.605 54.695 19.775 54.865 ;
        RECT 20.065 54.695 20.235 54.865 ;
        RECT 20.525 54.695 20.695 54.865 ;
        RECT 20.985 54.695 21.155 54.865 ;
        RECT 21.445 54.695 21.615 54.865 ;
        RECT 21.905 54.695 22.075 54.865 ;
        RECT 22.365 54.695 22.535 54.865 ;
        RECT 22.825 54.695 22.995 54.865 ;
        RECT 23.285 54.695 23.455 54.865 ;
        RECT 23.745 54.695 23.915 54.865 ;
        RECT 24.205 54.695 24.375 54.865 ;
        RECT 24.665 54.695 24.835 54.865 ;
        RECT 25.125 54.695 25.295 54.865 ;
        RECT 25.585 54.695 25.755 54.865 ;
        RECT 26.045 54.695 26.215 54.865 ;
        RECT 26.505 54.695 26.675 54.865 ;
        RECT 26.965 54.695 27.135 54.865 ;
        RECT 27.425 54.695 27.595 54.865 ;
        RECT 27.885 54.695 28.055 54.865 ;
        RECT 28.345 54.695 28.515 54.865 ;
        RECT 28.805 54.695 28.975 54.865 ;
        RECT 29.265 54.695 29.435 54.865 ;
        RECT 29.725 54.695 29.895 54.865 ;
        RECT 30.185 54.695 30.355 54.865 ;
        RECT 30.645 54.695 30.815 54.865 ;
        RECT 31.105 54.695 31.275 54.865 ;
        RECT 31.565 54.695 31.735 54.865 ;
        RECT 32.025 54.695 32.195 54.865 ;
        RECT 32.485 54.695 32.655 54.865 ;
        RECT 32.945 54.695 33.115 54.865 ;
        RECT 33.405 54.695 33.575 54.865 ;
        RECT 33.865 54.695 34.035 54.865 ;
        RECT 34.325 54.695 34.495 54.865 ;
        RECT 34.785 54.695 34.955 54.865 ;
        RECT 35.245 54.695 35.415 54.865 ;
        RECT 35.705 54.695 35.875 54.865 ;
        RECT 36.165 54.695 36.335 54.865 ;
        RECT 36.625 54.695 36.795 54.865 ;
        RECT 37.085 54.695 37.255 54.865 ;
        RECT 37.545 54.695 37.715 54.865 ;
        RECT 38.005 54.695 38.175 54.865 ;
        RECT 38.465 54.695 38.635 54.865 ;
        RECT 38.925 54.695 39.095 54.865 ;
        RECT 39.385 54.695 39.555 54.865 ;
        RECT 39.845 54.695 40.015 54.865 ;
        RECT 40.305 54.695 40.475 54.865 ;
        RECT 40.765 54.695 40.935 54.865 ;
        RECT 41.225 54.695 41.395 54.865 ;
        RECT 41.685 54.695 41.855 54.865 ;
        RECT 42.145 54.695 42.315 54.865 ;
        RECT 42.605 54.695 42.775 54.865 ;
        RECT 43.065 54.695 43.235 54.865 ;
        RECT 43.525 54.695 43.695 54.865 ;
        RECT 43.985 54.695 44.155 54.865 ;
        RECT 44.445 54.695 44.615 54.865 ;
        RECT 44.905 54.695 45.075 54.865 ;
        RECT 45.365 54.695 45.535 54.865 ;
        RECT 45.825 54.695 45.995 54.865 ;
        RECT 46.285 54.695 46.455 54.865 ;
        RECT 46.745 54.695 46.915 54.865 ;
        RECT 47.205 54.695 47.375 54.865 ;
        RECT 47.665 54.695 47.835 54.865 ;
        RECT 48.125 54.695 48.295 54.865 ;
        RECT 48.585 54.695 48.755 54.865 ;
        RECT 49.045 54.695 49.215 54.865 ;
        RECT 49.505 54.695 49.675 54.865 ;
        RECT 49.965 54.695 50.135 54.865 ;
        RECT 50.425 54.695 50.595 54.865 ;
        RECT 50.885 54.695 51.055 54.865 ;
        RECT 51.345 54.695 51.515 54.865 ;
        RECT 51.805 54.695 51.975 54.865 ;
        RECT 52.265 54.695 52.435 54.865 ;
        RECT 52.725 54.695 52.895 54.865 ;
        RECT 53.185 54.695 53.355 54.865 ;
        RECT 53.645 54.695 53.815 54.865 ;
        RECT 54.105 54.695 54.275 54.865 ;
        RECT 54.565 54.695 54.735 54.865 ;
        RECT 55.025 54.695 55.195 54.865 ;
        RECT 55.485 54.695 55.655 54.865 ;
        RECT 55.945 54.695 56.115 54.865 ;
        RECT 56.405 54.695 56.575 54.865 ;
        RECT 56.865 54.695 57.035 54.865 ;
        RECT 57.325 54.695 57.495 54.865 ;
        RECT 57.785 54.695 57.955 54.865 ;
        RECT 58.245 54.695 58.415 54.865 ;
        RECT 58.705 54.695 58.875 54.865 ;
        RECT 59.165 54.695 59.335 54.865 ;
        RECT 59.625 54.695 59.795 54.865 ;
        RECT 60.085 54.695 60.255 54.865 ;
        RECT 60.545 54.695 60.715 54.865 ;
        RECT 61.005 54.695 61.175 54.865 ;
        RECT 61.465 54.695 61.635 54.865 ;
        RECT 61.925 54.695 62.095 54.865 ;
        RECT 62.385 54.695 62.555 54.865 ;
        RECT 62.845 54.695 63.015 54.865 ;
        RECT 63.305 54.695 63.475 54.865 ;
        RECT 63.765 54.695 63.935 54.865 ;
        RECT 64.225 54.695 64.395 54.865 ;
        RECT 64.685 54.695 64.855 54.865 ;
        RECT 65.145 54.695 65.315 54.865 ;
        RECT 65.605 54.695 65.775 54.865 ;
        RECT 66.065 54.695 66.235 54.865 ;
        RECT 66.525 54.695 66.695 54.865 ;
        RECT 66.985 54.695 67.155 54.865 ;
        RECT 67.445 54.695 67.615 54.865 ;
        RECT 67.905 54.695 68.075 54.865 ;
        RECT 68.365 54.695 68.535 54.865 ;
        RECT 68.825 54.695 68.995 54.865 ;
        RECT 69.285 54.695 69.455 54.865 ;
        RECT 69.745 54.695 69.915 54.865 ;
        RECT 70.205 54.695 70.375 54.865 ;
        RECT 70.665 54.695 70.835 54.865 ;
        RECT 71.125 54.695 71.295 54.865 ;
        RECT 71.585 54.695 71.755 54.865 ;
        RECT 72.045 54.695 72.215 54.865 ;
        RECT 72.505 54.695 72.675 54.865 ;
        RECT 72.965 54.695 73.135 54.865 ;
        RECT 73.425 54.695 73.595 54.865 ;
        RECT 73.885 54.695 74.055 54.865 ;
        RECT 74.345 54.695 74.515 54.865 ;
        RECT 74.805 54.695 74.975 54.865 ;
        RECT 75.265 54.695 75.435 54.865 ;
        RECT 75.725 54.695 75.895 54.865 ;
        RECT 76.185 54.695 76.355 54.865 ;
        RECT 76.645 54.695 76.815 54.865 ;
        RECT 77.105 54.695 77.275 54.865 ;
        RECT 77.565 54.695 77.735 54.865 ;
        RECT 78.025 54.695 78.195 54.865 ;
        RECT 78.485 54.695 78.655 54.865 ;
        RECT 78.945 54.695 79.115 54.865 ;
        RECT 79.405 54.695 79.575 54.865 ;
        RECT 79.865 54.695 80.035 54.865 ;
        RECT 80.325 54.695 80.495 54.865 ;
        RECT 80.785 54.695 80.955 54.865 ;
        RECT 81.245 54.695 81.415 54.865 ;
        RECT 81.705 54.695 81.875 54.865 ;
        RECT 82.165 54.695 82.335 54.865 ;
        RECT 82.625 54.695 82.795 54.865 ;
        RECT 83.085 54.695 83.255 54.865 ;
        RECT 83.545 54.695 83.715 54.865 ;
        RECT 84.005 54.695 84.175 54.865 ;
        RECT 84.465 54.695 84.635 54.865 ;
        RECT 84.925 54.695 85.095 54.865 ;
        RECT 85.385 54.695 85.555 54.865 ;
        RECT 85.845 54.695 86.015 54.865 ;
        RECT 86.305 54.695 86.475 54.865 ;
        RECT 86.765 54.695 86.935 54.865 ;
        RECT 87.225 54.695 87.395 54.865 ;
        RECT 87.685 54.695 87.855 54.865 ;
        RECT 88.145 54.695 88.315 54.865 ;
        RECT 88.605 54.695 88.775 54.865 ;
        RECT 89.065 54.695 89.235 54.865 ;
        RECT 89.525 54.695 89.695 54.865 ;
        RECT 89.985 54.695 90.155 54.865 ;
        RECT 90.445 54.695 90.615 54.865 ;
        RECT 90.905 54.695 91.075 54.865 ;
        RECT 91.365 54.695 91.535 54.865 ;
        RECT 91.825 54.695 91.995 54.865 ;
        RECT 92.285 54.695 92.455 54.865 ;
        RECT 92.745 54.695 92.915 54.865 ;
        RECT 93.205 54.695 93.375 54.865 ;
        RECT 93.665 54.695 93.835 54.865 ;
        RECT 94.125 54.695 94.295 54.865 ;
        RECT 94.585 54.695 94.755 54.865 ;
        RECT 95.045 54.695 95.215 54.865 ;
        RECT 95.505 54.695 95.675 54.865 ;
        RECT 95.965 54.695 96.135 54.865 ;
        RECT 96.425 54.695 96.595 54.865 ;
        RECT 96.885 54.695 97.055 54.865 ;
        RECT 97.345 54.695 97.515 54.865 ;
        RECT 97.805 54.695 97.975 54.865 ;
        RECT 98.265 54.695 98.435 54.865 ;
        RECT 98.725 54.695 98.895 54.865 ;
        RECT 99.185 54.695 99.355 54.865 ;
        RECT 99.645 54.695 99.815 54.865 ;
        RECT 16.845 49.255 17.015 49.425 ;
        RECT 17.305 49.255 17.475 49.425 ;
        RECT 17.765 49.255 17.935 49.425 ;
        RECT 18.225 49.255 18.395 49.425 ;
        RECT 18.685 49.255 18.855 49.425 ;
        RECT 19.145 49.255 19.315 49.425 ;
        RECT 19.605 49.255 19.775 49.425 ;
        RECT 20.065 49.255 20.235 49.425 ;
        RECT 20.525 49.255 20.695 49.425 ;
        RECT 20.985 49.255 21.155 49.425 ;
        RECT 21.445 49.255 21.615 49.425 ;
        RECT 21.905 49.255 22.075 49.425 ;
        RECT 22.365 49.255 22.535 49.425 ;
        RECT 22.825 49.255 22.995 49.425 ;
        RECT 23.285 49.255 23.455 49.425 ;
        RECT 23.745 49.255 23.915 49.425 ;
        RECT 24.205 49.255 24.375 49.425 ;
        RECT 24.665 49.255 24.835 49.425 ;
        RECT 25.125 49.255 25.295 49.425 ;
        RECT 25.585 49.255 25.755 49.425 ;
        RECT 26.045 49.255 26.215 49.425 ;
        RECT 26.505 49.255 26.675 49.425 ;
        RECT 26.965 49.255 27.135 49.425 ;
        RECT 27.425 49.255 27.595 49.425 ;
        RECT 27.885 49.255 28.055 49.425 ;
        RECT 28.345 49.255 28.515 49.425 ;
        RECT 28.805 49.255 28.975 49.425 ;
        RECT 29.265 49.255 29.435 49.425 ;
        RECT 29.725 49.255 29.895 49.425 ;
        RECT 30.185 49.255 30.355 49.425 ;
        RECT 30.645 49.255 30.815 49.425 ;
        RECT 31.105 49.255 31.275 49.425 ;
        RECT 31.565 49.255 31.735 49.425 ;
        RECT 32.025 49.255 32.195 49.425 ;
        RECT 32.485 49.255 32.655 49.425 ;
        RECT 32.945 49.255 33.115 49.425 ;
        RECT 33.405 49.255 33.575 49.425 ;
        RECT 33.865 49.255 34.035 49.425 ;
        RECT 34.325 49.255 34.495 49.425 ;
        RECT 34.785 49.255 34.955 49.425 ;
        RECT 35.245 49.255 35.415 49.425 ;
        RECT 35.705 49.255 35.875 49.425 ;
        RECT 36.165 49.255 36.335 49.425 ;
        RECT 36.625 49.255 36.795 49.425 ;
        RECT 37.085 49.255 37.255 49.425 ;
        RECT 37.545 49.255 37.715 49.425 ;
        RECT 38.005 49.255 38.175 49.425 ;
        RECT 38.465 49.255 38.635 49.425 ;
        RECT 38.925 49.255 39.095 49.425 ;
        RECT 39.385 49.255 39.555 49.425 ;
        RECT 39.845 49.255 40.015 49.425 ;
        RECT 40.305 49.255 40.475 49.425 ;
        RECT 40.765 49.255 40.935 49.425 ;
        RECT 41.225 49.255 41.395 49.425 ;
        RECT 41.685 49.255 41.855 49.425 ;
        RECT 42.145 49.255 42.315 49.425 ;
        RECT 42.605 49.255 42.775 49.425 ;
        RECT 43.065 49.255 43.235 49.425 ;
        RECT 43.525 49.255 43.695 49.425 ;
        RECT 43.985 49.255 44.155 49.425 ;
        RECT 44.445 49.255 44.615 49.425 ;
        RECT 44.905 49.255 45.075 49.425 ;
        RECT 45.365 49.255 45.535 49.425 ;
        RECT 45.825 49.255 45.995 49.425 ;
        RECT 46.285 49.255 46.455 49.425 ;
        RECT 46.745 49.255 46.915 49.425 ;
        RECT 47.205 49.255 47.375 49.425 ;
        RECT 47.665 49.255 47.835 49.425 ;
        RECT 48.125 49.255 48.295 49.425 ;
        RECT 48.585 49.255 48.755 49.425 ;
        RECT 49.045 49.255 49.215 49.425 ;
        RECT 49.505 49.255 49.675 49.425 ;
        RECT 49.965 49.255 50.135 49.425 ;
        RECT 50.425 49.255 50.595 49.425 ;
        RECT 50.885 49.255 51.055 49.425 ;
        RECT 51.345 49.255 51.515 49.425 ;
        RECT 51.805 49.255 51.975 49.425 ;
        RECT 52.265 49.255 52.435 49.425 ;
        RECT 52.725 49.255 52.895 49.425 ;
        RECT 53.185 49.255 53.355 49.425 ;
        RECT 53.645 49.255 53.815 49.425 ;
        RECT 54.105 49.255 54.275 49.425 ;
        RECT 54.565 49.255 54.735 49.425 ;
        RECT 55.025 49.255 55.195 49.425 ;
        RECT 55.485 49.255 55.655 49.425 ;
        RECT 55.945 49.255 56.115 49.425 ;
        RECT 56.405 49.255 56.575 49.425 ;
        RECT 56.865 49.255 57.035 49.425 ;
        RECT 57.325 49.255 57.495 49.425 ;
        RECT 57.785 49.255 57.955 49.425 ;
        RECT 58.245 49.255 58.415 49.425 ;
        RECT 58.705 49.255 58.875 49.425 ;
        RECT 59.165 49.255 59.335 49.425 ;
        RECT 59.625 49.255 59.795 49.425 ;
        RECT 60.085 49.255 60.255 49.425 ;
        RECT 60.545 49.255 60.715 49.425 ;
        RECT 61.005 49.255 61.175 49.425 ;
        RECT 61.465 49.255 61.635 49.425 ;
        RECT 61.925 49.255 62.095 49.425 ;
        RECT 62.385 49.255 62.555 49.425 ;
        RECT 62.845 49.255 63.015 49.425 ;
        RECT 63.305 49.255 63.475 49.425 ;
        RECT 63.765 49.255 63.935 49.425 ;
        RECT 64.225 49.255 64.395 49.425 ;
        RECT 64.685 49.255 64.855 49.425 ;
        RECT 65.145 49.255 65.315 49.425 ;
        RECT 65.605 49.255 65.775 49.425 ;
        RECT 66.065 49.255 66.235 49.425 ;
        RECT 66.525 49.255 66.695 49.425 ;
        RECT 66.985 49.255 67.155 49.425 ;
        RECT 67.445 49.255 67.615 49.425 ;
        RECT 67.905 49.255 68.075 49.425 ;
        RECT 68.365 49.255 68.535 49.425 ;
        RECT 68.825 49.255 68.995 49.425 ;
        RECT 69.285 49.255 69.455 49.425 ;
        RECT 69.745 49.255 69.915 49.425 ;
        RECT 70.205 49.255 70.375 49.425 ;
        RECT 70.665 49.255 70.835 49.425 ;
        RECT 71.125 49.255 71.295 49.425 ;
        RECT 71.585 49.255 71.755 49.425 ;
        RECT 72.045 49.255 72.215 49.425 ;
        RECT 72.505 49.255 72.675 49.425 ;
        RECT 72.965 49.255 73.135 49.425 ;
        RECT 73.425 49.255 73.595 49.425 ;
        RECT 73.885 49.255 74.055 49.425 ;
        RECT 74.345 49.255 74.515 49.425 ;
        RECT 74.805 49.255 74.975 49.425 ;
        RECT 75.265 49.255 75.435 49.425 ;
        RECT 75.725 49.255 75.895 49.425 ;
        RECT 76.185 49.255 76.355 49.425 ;
        RECT 76.645 49.255 76.815 49.425 ;
        RECT 77.105 49.255 77.275 49.425 ;
        RECT 77.565 49.255 77.735 49.425 ;
        RECT 78.025 49.255 78.195 49.425 ;
        RECT 78.485 49.255 78.655 49.425 ;
        RECT 78.945 49.255 79.115 49.425 ;
        RECT 79.405 49.255 79.575 49.425 ;
        RECT 79.865 49.255 80.035 49.425 ;
        RECT 80.325 49.255 80.495 49.425 ;
        RECT 80.785 49.255 80.955 49.425 ;
        RECT 81.245 49.255 81.415 49.425 ;
        RECT 81.705 49.255 81.875 49.425 ;
        RECT 82.165 49.255 82.335 49.425 ;
        RECT 82.625 49.255 82.795 49.425 ;
        RECT 83.085 49.255 83.255 49.425 ;
        RECT 83.545 49.255 83.715 49.425 ;
        RECT 84.005 49.255 84.175 49.425 ;
        RECT 84.465 49.255 84.635 49.425 ;
        RECT 84.925 49.255 85.095 49.425 ;
        RECT 85.385 49.255 85.555 49.425 ;
        RECT 85.845 49.255 86.015 49.425 ;
        RECT 86.305 49.255 86.475 49.425 ;
        RECT 86.765 49.255 86.935 49.425 ;
        RECT 87.225 49.255 87.395 49.425 ;
        RECT 87.685 49.255 87.855 49.425 ;
        RECT 88.145 49.255 88.315 49.425 ;
        RECT 88.605 49.255 88.775 49.425 ;
        RECT 89.065 49.255 89.235 49.425 ;
        RECT 89.525 49.255 89.695 49.425 ;
        RECT 89.985 49.255 90.155 49.425 ;
        RECT 90.445 49.255 90.615 49.425 ;
        RECT 90.905 49.255 91.075 49.425 ;
        RECT 91.365 49.255 91.535 49.425 ;
        RECT 91.825 49.255 91.995 49.425 ;
        RECT 92.285 49.255 92.455 49.425 ;
        RECT 92.745 49.255 92.915 49.425 ;
        RECT 93.205 49.255 93.375 49.425 ;
        RECT 93.665 49.255 93.835 49.425 ;
        RECT 94.125 49.255 94.295 49.425 ;
        RECT 94.585 49.255 94.755 49.425 ;
        RECT 95.045 49.255 95.215 49.425 ;
        RECT 95.505 49.255 95.675 49.425 ;
        RECT 95.965 49.255 96.135 49.425 ;
        RECT 96.425 49.255 96.595 49.425 ;
        RECT 96.885 49.255 97.055 49.425 ;
        RECT 97.345 49.255 97.515 49.425 ;
        RECT 97.805 49.255 97.975 49.425 ;
        RECT 98.265 49.255 98.435 49.425 ;
        RECT 98.725 49.255 98.895 49.425 ;
        RECT 99.185 49.255 99.355 49.425 ;
        RECT 99.645 49.255 99.815 49.425 ;
        RECT 16.845 43.815 17.015 43.985 ;
        RECT 17.305 43.815 17.475 43.985 ;
        RECT 17.765 43.815 17.935 43.985 ;
        RECT 18.225 43.815 18.395 43.985 ;
        RECT 18.685 43.815 18.855 43.985 ;
        RECT 19.145 43.815 19.315 43.985 ;
        RECT 19.605 43.815 19.775 43.985 ;
        RECT 20.065 43.815 20.235 43.985 ;
        RECT 20.525 43.815 20.695 43.985 ;
        RECT 20.985 43.815 21.155 43.985 ;
        RECT 21.445 43.815 21.615 43.985 ;
        RECT 21.905 43.815 22.075 43.985 ;
        RECT 22.365 43.815 22.535 43.985 ;
        RECT 22.825 43.815 22.995 43.985 ;
        RECT 23.285 43.815 23.455 43.985 ;
        RECT 23.745 43.815 23.915 43.985 ;
        RECT 24.205 43.815 24.375 43.985 ;
        RECT 24.665 43.815 24.835 43.985 ;
        RECT 25.125 43.815 25.295 43.985 ;
        RECT 25.585 43.815 25.755 43.985 ;
        RECT 26.045 43.815 26.215 43.985 ;
        RECT 26.505 43.815 26.675 43.985 ;
        RECT 26.965 43.815 27.135 43.985 ;
        RECT 27.425 43.815 27.595 43.985 ;
        RECT 27.885 43.815 28.055 43.985 ;
        RECT 28.345 43.815 28.515 43.985 ;
        RECT 28.805 43.815 28.975 43.985 ;
        RECT 29.265 43.815 29.435 43.985 ;
        RECT 29.725 43.815 29.895 43.985 ;
        RECT 30.185 43.815 30.355 43.985 ;
        RECT 30.645 43.815 30.815 43.985 ;
        RECT 31.105 43.815 31.275 43.985 ;
        RECT 31.565 43.815 31.735 43.985 ;
        RECT 32.025 43.815 32.195 43.985 ;
        RECT 32.485 43.815 32.655 43.985 ;
        RECT 32.945 43.815 33.115 43.985 ;
        RECT 33.405 43.815 33.575 43.985 ;
        RECT 33.865 43.815 34.035 43.985 ;
        RECT 34.325 43.815 34.495 43.985 ;
        RECT 34.785 43.815 34.955 43.985 ;
        RECT 35.245 43.815 35.415 43.985 ;
        RECT 35.705 43.815 35.875 43.985 ;
        RECT 36.165 43.815 36.335 43.985 ;
        RECT 36.625 43.815 36.795 43.985 ;
        RECT 37.085 43.815 37.255 43.985 ;
        RECT 37.545 43.815 37.715 43.985 ;
        RECT 38.005 43.815 38.175 43.985 ;
        RECT 38.465 43.815 38.635 43.985 ;
        RECT 38.925 43.815 39.095 43.985 ;
        RECT 39.385 43.815 39.555 43.985 ;
        RECT 39.845 43.815 40.015 43.985 ;
        RECT 40.305 43.815 40.475 43.985 ;
        RECT 40.765 43.815 40.935 43.985 ;
        RECT 41.225 43.815 41.395 43.985 ;
        RECT 41.685 43.815 41.855 43.985 ;
        RECT 42.145 43.815 42.315 43.985 ;
        RECT 42.605 43.815 42.775 43.985 ;
        RECT 43.065 43.815 43.235 43.985 ;
        RECT 43.525 43.815 43.695 43.985 ;
        RECT 43.985 43.815 44.155 43.985 ;
        RECT 44.445 43.815 44.615 43.985 ;
        RECT 44.905 43.815 45.075 43.985 ;
        RECT 45.365 43.815 45.535 43.985 ;
        RECT 45.825 43.815 45.995 43.985 ;
        RECT 46.285 43.815 46.455 43.985 ;
        RECT 46.745 43.815 46.915 43.985 ;
        RECT 47.205 43.815 47.375 43.985 ;
        RECT 47.665 43.815 47.835 43.985 ;
        RECT 48.125 43.815 48.295 43.985 ;
        RECT 48.585 43.815 48.755 43.985 ;
        RECT 49.045 43.815 49.215 43.985 ;
        RECT 49.505 43.815 49.675 43.985 ;
        RECT 49.965 43.815 50.135 43.985 ;
        RECT 50.425 43.815 50.595 43.985 ;
        RECT 50.885 43.815 51.055 43.985 ;
        RECT 51.345 43.815 51.515 43.985 ;
        RECT 51.805 43.815 51.975 43.985 ;
        RECT 52.265 43.815 52.435 43.985 ;
        RECT 52.725 43.815 52.895 43.985 ;
        RECT 53.185 43.815 53.355 43.985 ;
        RECT 53.645 43.815 53.815 43.985 ;
        RECT 54.105 43.815 54.275 43.985 ;
        RECT 54.565 43.815 54.735 43.985 ;
        RECT 55.025 43.815 55.195 43.985 ;
        RECT 55.485 43.815 55.655 43.985 ;
        RECT 55.945 43.815 56.115 43.985 ;
        RECT 56.405 43.815 56.575 43.985 ;
        RECT 56.865 43.815 57.035 43.985 ;
        RECT 57.325 43.815 57.495 43.985 ;
        RECT 57.785 43.815 57.955 43.985 ;
        RECT 58.245 43.815 58.415 43.985 ;
        RECT 58.705 43.815 58.875 43.985 ;
        RECT 59.165 43.815 59.335 43.985 ;
        RECT 59.625 43.815 59.795 43.985 ;
        RECT 60.085 43.815 60.255 43.985 ;
        RECT 60.545 43.815 60.715 43.985 ;
        RECT 61.005 43.815 61.175 43.985 ;
        RECT 61.465 43.815 61.635 43.985 ;
        RECT 61.925 43.815 62.095 43.985 ;
        RECT 62.385 43.815 62.555 43.985 ;
        RECT 62.845 43.815 63.015 43.985 ;
        RECT 63.305 43.815 63.475 43.985 ;
        RECT 63.765 43.815 63.935 43.985 ;
        RECT 64.225 43.815 64.395 43.985 ;
        RECT 64.685 43.815 64.855 43.985 ;
        RECT 65.145 43.815 65.315 43.985 ;
        RECT 65.605 43.815 65.775 43.985 ;
        RECT 66.065 43.815 66.235 43.985 ;
        RECT 66.525 43.815 66.695 43.985 ;
        RECT 66.985 43.815 67.155 43.985 ;
        RECT 67.445 43.815 67.615 43.985 ;
        RECT 67.905 43.815 68.075 43.985 ;
        RECT 68.365 43.815 68.535 43.985 ;
        RECT 68.825 43.815 68.995 43.985 ;
        RECT 69.285 43.815 69.455 43.985 ;
        RECT 69.745 43.815 69.915 43.985 ;
        RECT 70.205 43.815 70.375 43.985 ;
        RECT 70.665 43.815 70.835 43.985 ;
        RECT 71.125 43.815 71.295 43.985 ;
        RECT 71.585 43.815 71.755 43.985 ;
        RECT 72.045 43.815 72.215 43.985 ;
        RECT 72.505 43.815 72.675 43.985 ;
        RECT 72.965 43.815 73.135 43.985 ;
        RECT 73.425 43.815 73.595 43.985 ;
        RECT 73.885 43.815 74.055 43.985 ;
        RECT 74.345 43.815 74.515 43.985 ;
        RECT 74.805 43.815 74.975 43.985 ;
        RECT 75.265 43.815 75.435 43.985 ;
        RECT 75.725 43.815 75.895 43.985 ;
        RECT 76.185 43.815 76.355 43.985 ;
        RECT 76.645 43.815 76.815 43.985 ;
        RECT 77.105 43.815 77.275 43.985 ;
        RECT 77.565 43.815 77.735 43.985 ;
        RECT 78.025 43.815 78.195 43.985 ;
        RECT 78.485 43.815 78.655 43.985 ;
        RECT 78.945 43.815 79.115 43.985 ;
        RECT 79.405 43.815 79.575 43.985 ;
        RECT 79.865 43.815 80.035 43.985 ;
        RECT 80.325 43.815 80.495 43.985 ;
        RECT 80.785 43.815 80.955 43.985 ;
        RECT 81.245 43.815 81.415 43.985 ;
        RECT 81.705 43.815 81.875 43.985 ;
        RECT 82.165 43.815 82.335 43.985 ;
        RECT 82.625 43.815 82.795 43.985 ;
        RECT 83.085 43.815 83.255 43.985 ;
        RECT 83.545 43.815 83.715 43.985 ;
        RECT 84.005 43.815 84.175 43.985 ;
        RECT 84.465 43.815 84.635 43.985 ;
        RECT 84.925 43.815 85.095 43.985 ;
        RECT 85.385 43.815 85.555 43.985 ;
        RECT 85.845 43.815 86.015 43.985 ;
        RECT 86.305 43.815 86.475 43.985 ;
        RECT 86.765 43.815 86.935 43.985 ;
        RECT 87.225 43.815 87.395 43.985 ;
        RECT 87.685 43.815 87.855 43.985 ;
        RECT 88.145 43.815 88.315 43.985 ;
        RECT 88.605 43.815 88.775 43.985 ;
        RECT 89.065 43.815 89.235 43.985 ;
        RECT 89.525 43.815 89.695 43.985 ;
        RECT 89.985 43.815 90.155 43.985 ;
        RECT 90.445 43.815 90.615 43.985 ;
        RECT 90.905 43.815 91.075 43.985 ;
        RECT 91.365 43.815 91.535 43.985 ;
        RECT 91.825 43.815 91.995 43.985 ;
        RECT 92.285 43.815 92.455 43.985 ;
        RECT 92.745 43.815 92.915 43.985 ;
        RECT 93.205 43.815 93.375 43.985 ;
        RECT 93.665 43.815 93.835 43.985 ;
        RECT 94.125 43.815 94.295 43.985 ;
        RECT 94.585 43.815 94.755 43.985 ;
        RECT 95.045 43.815 95.215 43.985 ;
        RECT 95.505 43.815 95.675 43.985 ;
        RECT 95.965 43.815 96.135 43.985 ;
        RECT 96.425 43.815 96.595 43.985 ;
        RECT 96.885 43.815 97.055 43.985 ;
        RECT 97.345 43.815 97.515 43.985 ;
        RECT 97.805 43.815 97.975 43.985 ;
        RECT 98.265 43.815 98.435 43.985 ;
        RECT 98.725 43.815 98.895 43.985 ;
        RECT 99.185 43.815 99.355 43.985 ;
        RECT 99.645 43.815 99.815 43.985 ;
        RECT 16.845 38.375 17.015 38.545 ;
        RECT 17.305 38.375 17.475 38.545 ;
        RECT 17.765 38.375 17.935 38.545 ;
        RECT 18.225 38.375 18.395 38.545 ;
        RECT 18.685 38.375 18.855 38.545 ;
        RECT 19.145 38.375 19.315 38.545 ;
        RECT 19.605 38.375 19.775 38.545 ;
        RECT 20.065 38.375 20.235 38.545 ;
        RECT 20.525 38.375 20.695 38.545 ;
        RECT 20.985 38.375 21.155 38.545 ;
        RECT 21.445 38.375 21.615 38.545 ;
        RECT 21.905 38.375 22.075 38.545 ;
        RECT 22.365 38.375 22.535 38.545 ;
        RECT 22.825 38.375 22.995 38.545 ;
        RECT 23.285 38.375 23.455 38.545 ;
        RECT 23.745 38.375 23.915 38.545 ;
        RECT 24.205 38.375 24.375 38.545 ;
        RECT 24.665 38.375 24.835 38.545 ;
        RECT 25.125 38.375 25.295 38.545 ;
        RECT 25.585 38.375 25.755 38.545 ;
        RECT 26.045 38.375 26.215 38.545 ;
        RECT 26.505 38.375 26.675 38.545 ;
        RECT 26.965 38.375 27.135 38.545 ;
        RECT 27.425 38.375 27.595 38.545 ;
        RECT 27.885 38.375 28.055 38.545 ;
        RECT 28.345 38.375 28.515 38.545 ;
        RECT 28.805 38.375 28.975 38.545 ;
        RECT 29.265 38.375 29.435 38.545 ;
        RECT 29.725 38.375 29.895 38.545 ;
        RECT 30.185 38.375 30.355 38.545 ;
        RECT 30.645 38.375 30.815 38.545 ;
        RECT 31.105 38.375 31.275 38.545 ;
        RECT 31.565 38.375 31.735 38.545 ;
        RECT 32.025 38.375 32.195 38.545 ;
        RECT 32.485 38.375 32.655 38.545 ;
        RECT 32.945 38.375 33.115 38.545 ;
        RECT 33.405 38.375 33.575 38.545 ;
        RECT 33.865 38.375 34.035 38.545 ;
        RECT 34.325 38.375 34.495 38.545 ;
        RECT 34.785 38.375 34.955 38.545 ;
        RECT 35.245 38.375 35.415 38.545 ;
        RECT 35.705 38.375 35.875 38.545 ;
        RECT 36.165 38.375 36.335 38.545 ;
        RECT 36.625 38.375 36.795 38.545 ;
        RECT 37.085 38.375 37.255 38.545 ;
        RECT 37.545 38.375 37.715 38.545 ;
        RECT 38.005 38.375 38.175 38.545 ;
        RECT 38.465 38.375 38.635 38.545 ;
        RECT 38.925 38.375 39.095 38.545 ;
        RECT 39.385 38.375 39.555 38.545 ;
        RECT 39.845 38.375 40.015 38.545 ;
        RECT 40.305 38.375 40.475 38.545 ;
        RECT 40.765 38.375 40.935 38.545 ;
        RECT 41.225 38.375 41.395 38.545 ;
        RECT 41.685 38.375 41.855 38.545 ;
        RECT 42.145 38.375 42.315 38.545 ;
        RECT 42.605 38.375 42.775 38.545 ;
        RECT 43.065 38.375 43.235 38.545 ;
        RECT 43.525 38.375 43.695 38.545 ;
        RECT 43.985 38.375 44.155 38.545 ;
        RECT 44.445 38.375 44.615 38.545 ;
        RECT 44.905 38.375 45.075 38.545 ;
        RECT 45.365 38.375 45.535 38.545 ;
        RECT 45.825 38.375 45.995 38.545 ;
        RECT 46.285 38.375 46.455 38.545 ;
        RECT 46.745 38.375 46.915 38.545 ;
        RECT 47.205 38.375 47.375 38.545 ;
        RECT 47.665 38.375 47.835 38.545 ;
        RECT 48.125 38.375 48.295 38.545 ;
        RECT 48.585 38.375 48.755 38.545 ;
        RECT 49.045 38.375 49.215 38.545 ;
        RECT 49.505 38.375 49.675 38.545 ;
        RECT 49.965 38.375 50.135 38.545 ;
        RECT 50.425 38.375 50.595 38.545 ;
        RECT 50.885 38.375 51.055 38.545 ;
        RECT 51.345 38.375 51.515 38.545 ;
        RECT 51.805 38.375 51.975 38.545 ;
        RECT 52.265 38.375 52.435 38.545 ;
        RECT 52.725 38.375 52.895 38.545 ;
        RECT 53.185 38.375 53.355 38.545 ;
        RECT 53.645 38.375 53.815 38.545 ;
        RECT 54.105 38.375 54.275 38.545 ;
        RECT 54.565 38.375 54.735 38.545 ;
        RECT 55.025 38.375 55.195 38.545 ;
        RECT 55.485 38.375 55.655 38.545 ;
        RECT 55.945 38.375 56.115 38.545 ;
        RECT 56.405 38.375 56.575 38.545 ;
        RECT 56.865 38.375 57.035 38.545 ;
        RECT 57.325 38.375 57.495 38.545 ;
        RECT 57.785 38.375 57.955 38.545 ;
        RECT 58.245 38.375 58.415 38.545 ;
        RECT 58.705 38.375 58.875 38.545 ;
        RECT 59.165 38.375 59.335 38.545 ;
        RECT 59.625 38.375 59.795 38.545 ;
        RECT 60.085 38.375 60.255 38.545 ;
        RECT 60.545 38.375 60.715 38.545 ;
        RECT 61.005 38.375 61.175 38.545 ;
        RECT 61.465 38.375 61.635 38.545 ;
        RECT 61.925 38.375 62.095 38.545 ;
        RECT 62.385 38.375 62.555 38.545 ;
        RECT 62.845 38.375 63.015 38.545 ;
        RECT 63.305 38.375 63.475 38.545 ;
        RECT 63.765 38.375 63.935 38.545 ;
        RECT 64.225 38.375 64.395 38.545 ;
        RECT 64.685 38.375 64.855 38.545 ;
        RECT 65.145 38.375 65.315 38.545 ;
        RECT 65.605 38.375 65.775 38.545 ;
        RECT 66.065 38.375 66.235 38.545 ;
        RECT 66.525 38.375 66.695 38.545 ;
        RECT 66.985 38.375 67.155 38.545 ;
        RECT 67.445 38.375 67.615 38.545 ;
        RECT 67.905 38.375 68.075 38.545 ;
        RECT 68.365 38.375 68.535 38.545 ;
        RECT 68.825 38.375 68.995 38.545 ;
        RECT 69.285 38.375 69.455 38.545 ;
        RECT 69.745 38.375 69.915 38.545 ;
        RECT 70.205 38.375 70.375 38.545 ;
        RECT 70.665 38.375 70.835 38.545 ;
        RECT 71.125 38.375 71.295 38.545 ;
        RECT 71.585 38.375 71.755 38.545 ;
        RECT 72.045 38.375 72.215 38.545 ;
        RECT 72.505 38.375 72.675 38.545 ;
        RECT 72.965 38.375 73.135 38.545 ;
        RECT 73.425 38.375 73.595 38.545 ;
        RECT 73.885 38.375 74.055 38.545 ;
        RECT 74.345 38.375 74.515 38.545 ;
        RECT 74.805 38.375 74.975 38.545 ;
        RECT 75.265 38.375 75.435 38.545 ;
        RECT 75.725 38.375 75.895 38.545 ;
        RECT 76.185 38.375 76.355 38.545 ;
        RECT 76.645 38.375 76.815 38.545 ;
        RECT 77.105 38.375 77.275 38.545 ;
        RECT 77.565 38.375 77.735 38.545 ;
        RECT 78.025 38.375 78.195 38.545 ;
        RECT 78.485 38.375 78.655 38.545 ;
        RECT 78.945 38.375 79.115 38.545 ;
        RECT 79.405 38.375 79.575 38.545 ;
        RECT 79.865 38.375 80.035 38.545 ;
        RECT 80.325 38.375 80.495 38.545 ;
        RECT 80.785 38.375 80.955 38.545 ;
        RECT 81.245 38.375 81.415 38.545 ;
        RECT 81.705 38.375 81.875 38.545 ;
        RECT 82.165 38.375 82.335 38.545 ;
        RECT 82.625 38.375 82.795 38.545 ;
        RECT 83.085 38.375 83.255 38.545 ;
        RECT 83.545 38.375 83.715 38.545 ;
        RECT 84.005 38.375 84.175 38.545 ;
        RECT 84.465 38.375 84.635 38.545 ;
        RECT 84.925 38.375 85.095 38.545 ;
        RECT 85.385 38.375 85.555 38.545 ;
        RECT 85.845 38.375 86.015 38.545 ;
        RECT 86.305 38.375 86.475 38.545 ;
        RECT 86.765 38.375 86.935 38.545 ;
        RECT 87.225 38.375 87.395 38.545 ;
        RECT 87.685 38.375 87.855 38.545 ;
        RECT 88.145 38.375 88.315 38.545 ;
        RECT 88.605 38.375 88.775 38.545 ;
        RECT 89.065 38.375 89.235 38.545 ;
        RECT 89.525 38.375 89.695 38.545 ;
        RECT 89.985 38.375 90.155 38.545 ;
        RECT 90.445 38.375 90.615 38.545 ;
        RECT 90.905 38.375 91.075 38.545 ;
        RECT 91.365 38.375 91.535 38.545 ;
        RECT 91.825 38.375 91.995 38.545 ;
        RECT 92.285 38.375 92.455 38.545 ;
        RECT 92.745 38.375 92.915 38.545 ;
        RECT 93.205 38.375 93.375 38.545 ;
        RECT 93.665 38.375 93.835 38.545 ;
        RECT 94.125 38.375 94.295 38.545 ;
        RECT 94.585 38.375 94.755 38.545 ;
        RECT 95.045 38.375 95.215 38.545 ;
        RECT 95.505 38.375 95.675 38.545 ;
        RECT 95.965 38.375 96.135 38.545 ;
        RECT 96.425 38.375 96.595 38.545 ;
        RECT 96.885 38.375 97.055 38.545 ;
        RECT 97.345 38.375 97.515 38.545 ;
        RECT 97.805 38.375 97.975 38.545 ;
        RECT 98.265 38.375 98.435 38.545 ;
        RECT 98.725 38.375 98.895 38.545 ;
        RECT 99.185 38.375 99.355 38.545 ;
        RECT 99.645 38.375 99.815 38.545 ;
        RECT 16.845 32.935 17.015 33.105 ;
        RECT 17.305 32.935 17.475 33.105 ;
        RECT 17.765 32.935 17.935 33.105 ;
        RECT 18.225 32.935 18.395 33.105 ;
        RECT 18.685 32.935 18.855 33.105 ;
        RECT 19.145 32.935 19.315 33.105 ;
        RECT 19.605 32.935 19.775 33.105 ;
        RECT 20.065 32.935 20.235 33.105 ;
        RECT 20.525 32.935 20.695 33.105 ;
        RECT 20.985 32.935 21.155 33.105 ;
        RECT 21.445 32.935 21.615 33.105 ;
        RECT 21.905 32.935 22.075 33.105 ;
        RECT 22.365 32.935 22.535 33.105 ;
        RECT 22.825 32.935 22.995 33.105 ;
        RECT 23.285 32.935 23.455 33.105 ;
        RECT 23.745 32.935 23.915 33.105 ;
        RECT 24.205 32.935 24.375 33.105 ;
        RECT 24.665 32.935 24.835 33.105 ;
        RECT 25.125 32.935 25.295 33.105 ;
        RECT 25.585 32.935 25.755 33.105 ;
        RECT 26.045 32.935 26.215 33.105 ;
        RECT 26.505 32.935 26.675 33.105 ;
        RECT 26.965 32.935 27.135 33.105 ;
        RECT 27.425 32.935 27.595 33.105 ;
        RECT 27.885 32.935 28.055 33.105 ;
        RECT 28.345 32.935 28.515 33.105 ;
        RECT 28.805 32.935 28.975 33.105 ;
        RECT 29.265 32.935 29.435 33.105 ;
        RECT 29.725 32.935 29.895 33.105 ;
        RECT 30.185 32.935 30.355 33.105 ;
        RECT 30.645 32.935 30.815 33.105 ;
        RECT 31.105 32.935 31.275 33.105 ;
        RECT 31.565 32.935 31.735 33.105 ;
        RECT 32.025 32.935 32.195 33.105 ;
        RECT 32.485 32.935 32.655 33.105 ;
        RECT 32.945 32.935 33.115 33.105 ;
        RECT 33.405 32.935 33.575 33.105 ;
        RECT 33.865 32.935 34.035 33.105 ;
        RECT 34.325 32.935 34.495 33.105 ;
        RECT 34.785 32.935 34.955 33.105 ;
        RECT 35.245 32.935 35.415 33.105 ;
        RECT 35.705 32.935 35.875 33.105 ;
        RECT 36.165 32.935 36.335 33.105 ;
        RECT 36.625 32.935 36.795 33.105 ;
        RECT 37.085 32.935 37.255 33.105 ;
        RECT 37.545 32.935 37.715 33.105 ;
        RECT 38.005 32.935 38.175 33.105 ;
        RECT 38.465 32.935 38.635 33.105 ;
        RECT 38.925 32.935 39.095 33.105 ;
        RECT 39.385 32.935 39.555 33.105 ;
        RECT 39.845 32.935 40.015 33.105 ;
        RECT 40.305 32.935 40.475 33.105 ;
        RECT 40.765 32.935 40.935 33.105 ;
        RECT 41.225 32.935 41.395 33.105 ;
        RECT 41.685 32.935 41.855 33.105 ;
        RECT 42.145 32.935 42.315 33.105 ;
        RECT 42.605 32.935 42.775 33.105 ;
        RECT 43.065 32.935 43.235 33.105 ;
        RECT 43.525 32.935 43.695 33.105 ;
        RECT 43.985 32.935 44.155 33.105 ;
        RECT 44.445 32.935 44.615 33.105 ;
        RECT 44.905 32.935 45.075 33.105 ;
        RECT 45.365 32.935 45.535 33.105 ;
        RECT 45.825 32.935 45.995 33.105 ;
        RECT 46.285 32.935 46.455 33.105 ;
        RECT 46.745 32.935 46.915 33.105 ;
        RECT 47.205 32.935 47.375 33.105 ;
        RECT 47.665 32.935 47.835 33.105 ;
        RECT 48.125 32.935 48.295 33.105 ;
        RECT 48.585 32.935 48.755 33.105 ;
        RECT 49.045 32.935 49.215 33.105 ;
        RECT 49.505 32.935 49.675 33.105 ;
        RECT 49.965 32.935 50.135 33.105 ;
        RECT 50.425 32.935 50.595 33.105 ;
        RECT 50.885 32.935 51.055 33.105 ;
        RECT 51.345 32.935 51.515 33.105 ;
        RECT 51.805 32.935 51.975 33.105 ;
        RECT 52.265 32.935 52.435 33.105 ;
        RECT 52.725 32.935 52.895 33.105 ;
        RECT 53.185 32.935 53.355 33.105 ;
        RECT 53.645 32.935 53.815 33.105 ;
        RECT 54.105 32.935 54.275 33.105 ;
        RECT 54.565 32.935 54.735 33.105 ;
        RECT 55.025 32.935 55.195 33.105 ;
        RECT 55.485 32.935 55.655 33.105 ;
        RECT 55.945 32.935 56.115 33.105 ;
        RECT 56.405 32.935 56.575 33.105 ;
        RECT 56.865 32.935 57.035 33.105 ;
        RECT 57.325 32.935 57.495 33.105 ;
        RECT 57.785 32.935 57.955 33.105 ;
        RECT 58.245 32.935 58.415 33.105 ;
        RECT 58.705 32.935 58.875 33.105 ;
        RECT 59.165 32.935 59.335 33.105 ;
        RECT 59.625 32.935 59.795 33.105 ;
        RECT 60.085 32.935 60.255 33.105 ;
        RECT 60.545 32.935 60.715 33.105 ;
        RECT 61.005 32.935 61.175 33.105 ;
        RECT 61.465 32.935 61.635 33.105 ;
        RECT 61.925 32.935 62.095 33.105 ;
        RECT 62.385 32.935 62.555 33.105 ;
        RECT 62.845 32.935 63.015 33.105 ;
        RECT 63.305 32.935 63.475 33.105 ;
        RECT 63.765 32.935 63.935 33.105 ;
        RECT 64.225 32.935 64.395 33.105 ;
        RECT 64.685 32.935 64.855 33.105 ;
        RECT 65.145 32.935 65.315 33.105 ;
        RECT 65.605 32.935 65.775 33.105 ;
        RECT 66.065 32.935 66.235 33.105 ;
        RECT 66.525 32.935 66.695 33.105 ;
        RECT 66.985 32.935 67.155 33.105 ;
        RECT 67.445 32.935 67.615 33.105 ;
        RECT 67.905 32.935 68.075 33.105 ;
        RECT 68.365 32.935 68.535 33.105 ;
        RECT 68.825 32.935 68.995 33.105 ;
        RECT 69.285 32.935 69.455 33.105 ;
        RECT 69.745 32.935 69.915 33.105 ;
        RECT 70.205 32.935 70.375 33.105 ;
        RECT 70.665 32.935 70.835 33.105 ;
        RECT 71.125 32.935 71.295 33.105 ;
        RECT 71.585 32.935 71.755 33.105 ;
        RECT 72.045 32.935 72.215 33.105 ;
        RECT 72.505 32.935 72.675 33.105 ;
        RECT 72.965 32.935 73.135 33.105 ;
        RECT 73.425 32.935 73.595 33.105 ;
        RECT 73.885 32.935 74.055 33.105 ;
        RECT 74.345 32.935 74.515 33.105 ;
        RECT 74.805 32.935 74.975 33.105 ;
        RECT 75.265 32.935 75.435 33.105 ;
        RECT 75.725 32.935 75.895 33.105 ;
        RECT 76.185 32.935 76.355 33.105 ;
        RECT 76.645 32.935 76.815 33.105 ;
        RECT 77.105 32.935 77.275 33.105 ;
        RECT 77.565 32.935 77.735 33.105 ;
        RECT 78.025 32.935 78.195 33.105 ;
        RECT 78.485 32.935 78.655 33.105 ;
        RECT 78.945 32.935 79.115 33.105 ;
        RECT 79.405 32.935 79.575 33.105 ;
        RECT 79.865 32.935 80.035 33.105 ;
        RECT 80.325 32.935 80.495 33.105 ;
        RECT 80.785 32.935 80.955 33.105 ;
        RECT 81.245 32.935 81.415 33.105 ;
        RECT 81.705 32.935 81.875 33.105 ;
        RECT 82.165 32.935 82.335 33.105 ;
        RECT 82.625 32.935 82.795 33.105 ;
        RECT 83.085 32.935 83.255 33.105 ;
        RECT 83.545 32.935 83.715 33.105 ;
        RECT 84.005 32.935 84.175 33.105 ;
        RECT 84.465 32.935 84.635 33.105 ;
        RECT 84.925 32.935 85.095 33.105 ;
        RECT 85.385 32.935 85.555 33.105 ;
        RECT 85.845 32.935 86.015 33.105 ;
        RECT 86.305 32.935 86.475 33.105 ;
        RECT 86.765 32.935 86.935 33.105 ;
        RECT 87.225 32.935 87.395 33.105 ;
        RECT 87.685 32.935 87.855 33.105 ;
        RECT 88.145 32.935 88.315 33.105 ;
        RECT 88.605 32.935 88.775 33.105 ;
        RECT 89.065 32.935 89.235 33.105 ;
        RECT 89.525 32.935 89.695 33.105 ;
        RECT 89.985 32.935 90.155 33.105 ;
        RECT 90.445 32.935 90.615 33.105 ;
        RECT 90.905 32.935 91.075 33.105 ;
        RECT 91.365 32.935 91.535 33.105 ;
        RECT 91.825 32.935 91.995 33.105 ;
        RECT 92.285 32.935 92.455 33.105 ;
        RECT 92.745 32.935 92.915 33.105 ;
        RECT 93.205 32.935 93.375 33.105 ;
        RECT 93.665 32.935 93.835 33.105 ;
        RECT 94.125 32.935 94.295 33.105 ;
        RECT 94.585 32.935 94.755 33.105 ;
        RECT 95.045 32.935 95.215 33.105 ;
        RECT 95.505 32.935 95.675 33.105 ;
        RECT 95.965 32.935 96.135 33.105 ;
        RECT 96.425 32.935 96.595 33.105 ;
        RECT 96.885 32.935 97.055 33.105 ;
        RECT 97.345 32.935 97.515 33.105 ;
        RECT 97.805 32.935 97.975 33.105 ;
        RECT 98.265 32.935 98.435 33.105 ;
        RECT 98.725 32.935 98.895 33.105 ;
        RECT 99.185 32.935 99.355 33.105 ;
        RECT 99.645 32.935 99.815 33.105 ;
        RECT 16.845 27.495 17.015 27.665 ;
        RECT 17.305 27.495 17.475 27.665 ;
        RECT 17.765 27.495 17.935 27.665 ;
        RECT 18.225 27.495 18.395 27.665 ;
        RECT 18.685 27.495 18.855 27.665 ;
        RECT 19.145 27.495 19.315 27.665 ;
        RECT 19.605 27.495 19.775 27.665 ;
        RECT 20.065 27.495 20.235 27.665 ;
        RECT 20.525 27.495 20.695 27.665 ;
        RECT 20.985 27.495 21.155 27.665 ;
        RECT 21.445 27.495 21.615 27.665 ;
        RECT 21.905 27.495 22.075 27.665 ;
        RECT 22.365 27.495 22.535 27.665 ;
        RECT 22.825 27.495 22.995 27.665 ;
        RECT 23.285 27.495 23.455 27.665 ;
        RECT 23.745 27.495 23.915 27.665 ;
        RECT 24.205 27.495 24.375 27.665 ;
        RECT 24.665 27.495 24.835 27.665 ;
        RECT 25.125 27.495 25.295 27.665 ;
        RECT 25.585 27.495 25.755 27.665 ;
        RECT 26.045 27.495 26.215 27.665 ;
        RECT 26.505 27.495 26.675 27.665 ;
        RECT 26.965 27.495 27.135 27.665 ;
        RECT 27.425 27.495 27.595 27.665 ;
        RECT 27.885 27.495 28.055 27.665 ;
        RECT 28.345 27.495 28.515 27.665 ;
        RECT 28.805 27.495 28.975 27.665 ;
        RECT 29.265 27.495 29.435 27.665 ;
        RECT 29.725 27.495 29.895 27.665 ;
        RECT 30.185 27.495 30.355 27.665 ;
        RECT 30.645 27.495 30.815 27.665 ;
        RECT 31.105 27.495 31.275 27.665 ;
        RECT 31.565 27.495 31.735 27.665 ;
        RECT 32.025 27.495 32.195 27.665 ;
        RECT 32.485 27.495 32.655 27.665 ;
        RECT 32.945 27.495 33.115 27.665 ;
        RECT 33.405 27.495 33.575 27.665 ;
        RECT 33.865 27.495 34.035 27.665 ;
        RECT 34.325 27.495 34.495 27.665 ;
        RECT 34.785 27.495 34.955 27.665 ;
        RECT 35.245 27.495 35.415 27.665 ;
        RECT 35.705 27.495 35.875 27.665 ;
        RECT 36.165 27.495 36.335 27.665 ;
        RECT 36.625 27.495 36.795 27.665 ;
        RECT 37.085 27.495 37.255 27.665 ;
        RECT 37.545 27.495 37.715 27.665 ;
        RECT 38.005 27.495 38.175 27.665 ;
        RECT 38.465 27.495 38.635 27.665 ;
        RECT 38.925 27.495 39.095 27.665 ;
        RECT 39.385 27.495 39.555 27.665 ;
        RECT 39.845 27.495 40.015 27.665 ;
        RECT 40.305 27.495 40.475 27.665 ;
        RECT 40.765 27.495 40.935 27.665 ;
        RECT 41.225 27.495 41.395 27.665 ;
        RECT 41.685 27.495 41.855 27.665 ;
        RECT 42.145 27.495 42.315 27.665 ;
        RECT 42.605 27.495 42.775 27.665 ;
        RECT 43.065 27.495 43.235 27.665 ;
        RECT 43.525 27.495 43.695 27.665 ;
        RECT 43.985 27.495 44.155 27.665 ;
        RECT 44.445 27.495 44.615 27.665 ;
        RECT 44.905 27.495 45.075 27.665 ;
        RECT 45.365 27.495 45.535 27.665 ;
        RECT 45.825 27.495 45.995 27.665 ;
        RECT 46.285 27.495 46.455 27.665 ;
        RECT 46.745 27.495 46.915 27.665 ;
        RECT 47.205 27.495 47.375 27.665 ;
        RECT 47.665 27.495 47.835 27.665 ;
        RECT 48.125 27.495 48.295 27.665 ;
        RECT 48.585 27.495 48.755 27.665 ;
        RECT 49.045 27.495 49.215 27.665 ;
        RECT 49.505 27.495 49.675 27.665 ;
        RECT 49.965 27.495 50.135 27.665 ;
        RECT 50.425 27.495 50.595 27.665 ;
        RECT 50.885 27.495 51.055 27.665 ;
        RECT 51.345 27.495 51.515 27.665 ;
        RECT 51.805 27.495 51.975 27.665 ;
        RECT 52.265 27.495 52.435 27.665 ;
        RECT 52.725 27.495 52.895 27.665 ;
        RECT 53.185 27.495 53.355 27.665 ;
        RECT 53.645 27.495 53.815 27.665 ;
        RECT 54.105 27.495 54.275 27.665 ;
        RECT 54.565 27.495 54.735 27.665 ;
        RECT 55.025 27.495 55.195 27.665 ;
        RECT 55.485 27.495 55.655 27.665 ;
        RECT 55.945 27.495 56.115 27.665 ;
        RECT 56.405 27.495 56.575 27.665 ;
        RECT 56.865 27.495 57.035 27.665 ;
        RECT 57.325 27.495 57.495 27.665 ;
        RECT 57.785 27.495 57.955 27.665 ;
        RECT 58.245 27.495 58.415 27.665 ;
        RECT 58.705 27.495 58.875 27.665 ;
        RECT 59.165 27.495 59.335 27.665 ;
        RECT 59.625 27.495 59.795 27.665 ;
        RECT 60.085 27.495 60.255 27.665 ;
        RECT 60.545 27.495 60.715 27.665 ;
        RECT 61.005 27.495 61.175 27.665 ;
        RECT 61.465 27.495 61.635 27.665 ;
        RECT 61.925 27.495 62.095 27.665 ;
        RECT 62.385 27.495 62.555 27.665 ;
        RECT 62.845 27.495 63.015 27.665 ;
        RECT 63.305 27.495 63.475 27.665 ;
        RECT 63.765 27.495 63.935 27.665 ;
        RECT 64.225 27.495 64.395 27.665 ;
        RECT 64.685 27.495 64.855 27.665 ;
        RECT 65.145 27.495 65.315 27.665 ;
        RECT 65.605 27.495 65.775 27.665 ;
        RECT 66.065 27.495 66.235 27.665 ;
        RECT 66.525 27.495 66.695 27.665 ;
        RECT 66.985 27.495 67.155 27.665 ;
        RECT 67.445 27.495 67.615 27.665 ;
        RECT 67.905 27.495 68.075 27.665 ;
        RECT 68.365 27.495 68.535 27.665 ;
        RECT 68.825 27.495 68.995 27.665 ;
        RECT 69.285 27.495 69.455 27.665 ;
        RECT 69.745 27.495 69.915 27.665 ;
        RECT 70.205 27.495 70.375 27.665 ;
        RECT 70.665 27.495 70.835 27.665 ;
        RECT 71.125 27.495 71.295 27.665 ;
        RECT 71.585 27.495 71.755 27.665 ;
        RECT 72.045 27.495 72.215 27.665 ;
        RECT 72.505 27.495 72.675 27.665 ;
        RECT 72.965 27.495 73.135 27.665 ;
        RECT 73.425 27.495 73.595 27.665 ;
        RECT 73.885 27.495 74.055 27.665 ;
        RECT 74.345 27.495 74.515 27.665 ;
        RECT 74.805 27.495 74.975 27.665 ;
        RECT 75.265 27.495 75.435 27.665 ;
        RECT 75.725 27.495 75.895 27.665 ;
        RECT 76.185 27.495 76.355 27.665 ;
        RECT 76.645 27.495 76.815 27.665 ;
        RECT 77.105 27.495 77.275 27.665 ;
        RECT 77.565 27.495 77.735 27.665 ;
        RECT 78.025 27.495 78.195 27.665 ;
        RECT 78.485 27.495 78.655 27.665 ;
        RECT 78.945 27.495 79.115 27.665 ;
        RECT 79.405 27.495 79.575 27.665 ;
        RECT 79.865 27.495 80.035 27.665 ;
        RECT 80.325 27.495 80.495 27.665 ;
        RECT 80.785 27.495 80.955 27.665 ;
        RECT 81.245 27.495 81.415 27.665 ;
        RECT 81.705 27.495 81.875 27.665 ;
        RECT 82.165 27.495 82.335 27.665 ;
        RECT 82.625 27.495 82.795 27.665 ;
        RECT 83.085 27.495 83.255 27.665 ;
        RECT 83.545 27.495 83.715 27.665 ;
        RECT 84.005 27.495 84.175 27.665 ;
        RECT 84.465 27.495 84.635 27.665 ;
        RECT 84.925 27.495 85.095 27.665 ;
        RECT 85.385 27.495 85.555 27.665 ;
        RECT 85.845 27.495 86.015 27.665 ;
        RECT 86.305 27.495 86.475 27.665 ;
        RECT 86.765 27.495 86.935 27.665 ;
        RECT 87.225 27.495 87.395 27.665 ;
        RECT 87.685 27.495 87.855 27.665 ;
        RECT 88.145 27.495 88.315 27.665 ;
        RECT 88.605 27.495 88.775 27.665 ;
        RECT 89.065 27.495 89.235 27.665 ;
        RECT 89.525 27.495 89.695 27.665 ;
        RECT 89.985 27.495 90.155 27.665 ;
        RECT 90.445 27.495 90.615 27.665 ;
        RECT 90.905 27.495 91.075 27.665 ;
        RECT 91.365 27.495 91.535 27.665 ;
        RECT 91.825 27.495 91.995 27.665 ;
        RECT 92.285 27.495 92.455 27.665 ;
        RECT 92.745 27.495 92.915 27.665 ;
        RECT 93.205 27.495 93.375 27.665 ;
        RECT 93.665 27.495 93.835 27.665 ;
        RECT 94.125 27.495 94.295 27.665 ;
        RECT 94.585 27.495 94.755 27.665 ;
        RECT 95.045 27.495 95.215 27.665 ;
        RECT 95.505 27.495 95.675 27.665 ;
        RECT 95.965 27.495 96.135 27.665 ;
        RECT 96.425 27.495 96.595 27.665 ;
        RECT 96.885 27.495 97.055 27.665 ;
        RECT 97.345 27.495 97.515 27.665 ;
        RECT 97.805 27.495 97.975 27.665 ;
        RECT 98.265 27.495 98.435 27.665 ;
        RECT 98.725 27.495 98.895 27.665 ;
        RECT 99.185 27.495 99.355 27.665 ;
        RECT 99.645 27.495 99.815 27.665 ;
        RECT 16.845 22.055 17.015 22.225 ;
        RECT 17.305 22.055 17.475 22.225 ;
        RECT 17.765 22.055 17.935 22.225 ;
        RECT 18.225 22.055 18.395 22.225 ;
        RECT 18.685 22.055 18.855 22.225 ;
        RECT 19.145 22.055 19.315 22.225 ;
        RECT 19.605 22.055 19.775 22.225 ;
        RECT 20.065 22.055 20.235 22.225 ;
        RECT 20.525 22.055 20.695 22.225 ;
        RECT 20.985 22.055 21.155 22.225 ;
        RECT 21.445 22.055 21.615 22.225 ;
        RECT 21.905 22.055 22.075 22.225 ;
        RECT 22.365 22.055 22.535 22.225 ;
        RECT 22.825 22.055 22.995 22.225 ;
        RECT 23.285 22.055 23.455 22.225 ;
        RECT 23.745 22.055 23.915 22.225 ;
        RECT 24.205 22.055 24.375 22.225 ;
        RECT 24.665 22.055 24.835 22.225 ;
        RECT 25.125 22.055 25.295 22.225 ;
        RECT 25.585 22.055 25.755 22.225 ;
        RECT 26.045 22.055 26.215 22.225 ;
        RECT 26.505 22.055 26.675 22.225 ;
        RECT 26.965 22.055 27.135 22.225 ;
        RECT 27.425 22.055 27.595 22.225 ;
        RECT 27.885 22.055 28.055 22.225 ;
        RECT 28.345 22.055 28.515 22.225 ;
        RECT 28.805 22.055 28.975 22.225 ;
        RECT 29.265 22.055 29.435 22.225 ;
        RECT 29.725 22.055 29.895 22.225 ;
        RECT 30.185 22.055 30.355 22.225 ;
        RECT 30.645 22.055 30.815 22.225 ;
        RECT 31.105 22.055 31.275 22.225 ;
        RECT 31.565 22.055 31.735 22.225 ;
        RECT 32.025 22.055 32.195 22.225 ;
        RECT 32.485 22.055 32.655 22.225 ;
        RECT 32.945 22.055 33.115 22.225 ;
        RECT 33.405 22.055 33.575 22.225 ;
        RECT 33.865 22.055 34.035 22.225 ;
        RECT 34.325 22.055 34.495 22.225 ;
        RECT 34.785 22.055 34.955 22.225 ;
        RECT 35.245 22.055 35.415 22.225 ;
        RECT 35.705 22.055 35.875 22.225 ;
        RECT 36.165 22.055 36.335 22.225 ;
        RECT 36.625 22.055 36.795 22.225 ;
        RECT 37.085 22.055 37.255 22.225 ;
        RECT 37.545 22.055 37.715 22.225 ;
        RECT 38.005 22.055 38.175 22.225 ;
        RECT 38.465 22.055 38.635 22.225 ;
        RECT 38.925 22.055 39.095 22.225 ;
        RECT 39.385 22.055 39.555 22.225 ;
        RECT 39.845 22.055 40.015 22.225 ;
        RECT 40.305 22.055 40.475 22.225 ;
        RECT 40.765 22.055 40.935 22.225 ;
        RECT 41.225 22.055 41.395 22.225 ;
        RECT 41.685 22.055 41.855 22.225 ;
        RECT 42.145 22.055 42.315 22.225 ;
        RECT 42.605 22.055 42.775 22.225 ;
        RECT 43.065 22.055 43.235 22.225 ;
        RECT 43.525 22.055 43.695 22.225 ;
        RECT 43.985 22.055 44.155 22.225 ;
        RECT 44.445 22.055 44.615 22.225 ;
        RECT 44.905 22.055 45.075 22.225 ;
        RECT 45.365 22.055 45.535 22.225 ;
        RECT 45.825 22.055 45.995 22.225 ;
        RECT 46.285 22.055 46.455 22.225 ;
        RECT 46.745 22.055 46.915 22.225 ;
        RECT 47.205 22.055 47.375 22.225 ;
        RECT 47.665 22.055 47.835 22.225 ;
        RECT 48.125 22.055 48.295 22.225 ;
        RECT 48.585 22.055 48.755 22.225 ;
        RECT 49.045 22.055 49.215 22.225 ;
        RECT 49.505 22.055 49.675 22.225 ;
        RECT 49.965 22.055 50.135 22.225 ;
        RECT 50.425 22.055 50.595 22.225 ;
        RECT 50.885 22.055 51.055 22.225 ;
        RECT 51.345 22.055 51.515 22.225 ;
        RECT 51.805 22.055 51.975 22.225 ;
        RECT 52.265 22.055 52.435 22.225 ;
        RECT 52.725 22.055 52.895 22.225 ;
        RECT 53.185 22.055 53.355 22.225 ;
        RECT 53.645 22.055 53.815 22.225 ;
        RECT 54.105 22.055 54.275 22.225 ;
        RECT 54.565 22.055 54.735 22.225 ;
        RECT 55.025 22.055 55.195 22.225 ;
        RECT 55.485 22.055 55.655 22.225 ;
        RECT 55.945 22.055 56.115 22.225 ;
        RECT 56.405 22.055 56.575 22.225 ;
        RECT 56.865 22.055 57.035 22.225 ;
        RECT 57.325 22.055 57.495 22.225 ;
        RECT 57.785 22.055 57.955 22.225 ;
        RECT 58.245 22.055 58.415 22.225 ;
        RECT 58.705 22.055 58.875 22.225 ;
        RECT 59.165 22.055 59.335 22.225 ;
        RECT 59.625 22.055 59.795 22.225 ;
        RECT 60.085 22.055 60.255 22.225 ;
        RECT 60.545 22.055 60.715 22.225 ;
        RECT 61.005 22.055 61.175 22.225 ;
        RECT 61.465 22.055 61.635 22.225 ;
        RECT 61.925 22.055 62.095 22.225 ;
        RECT 62.385 22.055 62.555 22.225 ;
        RECT 62.845 22.055 63.015 22.225 ;
        RECT 63.305 22.055 63.475 22.225 ;
        RECT 63.765 22.055 63.935 22.225 ;
        RECT 64.225 22.055 64.395 22.225 ;
        RECT 64.685 22.055 64.855 22.225 ;
        RECT 65.145 22.055 65.315 22.225 ;
        RECT 65.605 22.055 65.775 22.225 ;
        RECT 66.065 22.055 66.235 22.225 ;
        RECT 66.525 22.055 66.695 22.225 ;
        RECT 66.985 22.055 67.155 22.225 ;
        RECT 67.445 22.055 67.615 22.225 ;
        RECT 67.905 22.055 68.075 22.225 ;
        RECT 68.365 22.055 68.535 22.225 ;
        RECT 68.825 22.055 68.995 22.225 ;
        RECT 69.285 22.055 69.455 22.225 ;
        RECT 69.745 22.055 69.915 22.225 ;
        RECT 70.205 22.055 70.375 22.225 ;
        RECT 70.665 22.055 70.835 22.225 ;
        RECT 71.125 22.055 71.295 22.225 ;
        RECT 71.585 22.055 71.755 22.225 ;
        RECT 72.045 22.055 72.215 22.225 ;
        RECT 72.505 22.055 72.675 22.225 ;
        RECT 72.965 22.055 73.135 22.225 ;
        RECT 73.425 22.055 73.595 22.225 ;
        RECT 73.885 22.055 74.055 22.225 ;
        RECT 74.345 22.055 74.515 22.225 ;
        RECT 74.805 22.055 74.975 22.225 ;
        RECT 75.265 22.055 75.435 22.225 ;
        RECT 75.725 22.055 75.895 22.225 ;
        RECT 76.185 22.055 76.355 22.225 ;
        RECT 76.645 22.055 76.815 22.225 ;
        RECT 77.105 22.055 77.275 22.225 ;
        RECT 77.565 22.055 77.735 22.225 ;
        RECT 78.025 22.055 78.195 22.225 ;
        RECT 78.485 22.055 78.655 22.225 ;
        RECT 78.945 22.055 79.115 22.225 ;
        RECT 79.405 22.055 79.575 22.225 ;
        RECT 79.865 22.055 80.035 22.225 ;
        RECT 80.325 22.055 80.495 22.225 ;
        RECT 80.785 22.055 80.955 22.225 ;
        RECT 81.245 22.055 81.415 22.225 ;
        RECT 81.705 22.055 81.875 22.225 ;
        RECT 82.165 22.055 82.335 22.225 ;
        RECT 82.625 22.055 82.795 22.225 ;
        RECT 83.085 22.055 83.255 22.225 ;
        RECT 83.545 22.055 83.715 22.225 ;
        RECT 84.005 22.055 84.175 22.225 ;
        RECT 84.465 22.055 84.635 22.225 ;
        RECT 84.925 22.055 85.095 22.225 ;
        RECT 85.385 22.055 85.555 22.225 ;
        RECT 85.845 22.055 86.015 22.225 ;
        RECT 86.305 22.055 86.475 22.225 ;
        RECT 86.765 22.055 86.935 22.225 ;
        RECT 87.225 22.055 87.395 22.225 ;
        RECT 87.685 22.055 87.855 22.225 ;
        RECT 88.145 22.055 88.315 22.225 ;
        RECT 88.605 22.055 88.775 22.225 ;
        RECT 89.065 22.055 89.235 22.225 ;
        RECT 89.525 22.055 89.695 22.225 ;
        RECT 89.985 22.055 90.155 22.225 ;
        RECT 90.445 22.055 90.615 22.225 ;
        RECT 90.905 22.055 91.075 22.225 ;
        RECT 91.365 22.055 91.535 22.225 ;
        RECT 91.825 22.055 91.995 22.225 ;
        RECT 92.285 22.055 92.455 22.225 ;
        RECT 92.745 22.055 92.915 22.225 ;
        RECT 93.205 22.055 93.375 22.225 ;
        RECT 93.665 22.055 93.835 22.225 ;
        RECT 94.125 22.055 94.295 22.225 ;
        RECT 94.585 22.055 94.755 22.225 ;
        RECT 95.045 22.055 95.215 22.225 ;
        RECT 95.505 22.055 95.675 22.225 ;
        RECT 95.965 22.055 96.135 22.225 ;
        RECT 96.425 22.055 96.595 22.225 ;
        RECT 96.885 22.055 97.055 22.225 ;
        RECT 97.345 22.055 97.515 22.225 ;
        RECT 97.805 22.055 97.975 22.225 ;
        RECT 98.265 22.055 98.435 22.225 ;
        RECT 98.725 22.055 98.895 22.225 ;
        RECT 99.185 22.055 99.355 22.225 ;
        RECT 99.645 22.055 99.815 22.225 ;
        RECT 16.845 16.615 17.015 16.785 ;
        RECT 17.305 16.615 17.475 16.785 ;
        RECT 17.765 16.615 17.935 16.785 ;
        RECT 18.225 16.615 18.395 16.785 ;
        RECT 18.685 16.615 18.855 16.785 ;
        RECT 19.145 16.615 19.315 16.785 ;
        RECT 19.605 16.615 19.775 16.785 ;
        RECT 20.065 16.615 20.235 16.785 ;
        RECT 20.525 16.615 20.695 16.785 ;
        RECT 20.985 16.615 21.155 16.785 ;
        RECT 21.445 16.615 21.615 16.785 ;
        RECT 21.905 16.615 22.075 16.785 ;
        RECT 22.365 16.615 22.535 16.785 ;
        RECT 22.825 16.615 22.995 16.785 ;
        RECT 23.285 16.615 23.455 16.785 ;
        RECT 23.745 16.615 23.915 16.785 ;
        RECT 24.205 16.615 24.375 16.785 ;
        RECT 24.665 16.615 24.835 16.785 ;
        RECT 25.125 16.615 25.295 16.785 ;
        RECT 25.585 16.615 25.755 16.785 ;
        RECT 26.045 16.615 26.215 16.785 ;
        RECT 26.505 16.615 26.675 16.785 ;
        RECT 26.965 16.615 27.135 16.785 ;
        RECT 27.425 16.615 27.595 16.785 ;
        RECT 27.885 16.615 28.055 16.785 ;
        RECT 28.345 16.615 28.515 16.785 ;
        RECT 28.805 16.615 28.975 16.785 ;
        RECT 29.265 16.615 29.435 16.785 ;
        RECT 29.725 16.615 29.895 16.785 ;
        RECT 30.185 16.615 30.355 16.785 ;
        RECT 30.645 16.615 30.815 16.785 ;
        RECT 31.105 16.615 31.275 16.785 ;
        RECT 31.565 16.615 31.735 16.785 ;
        RECT 32.025 16.615 32.195 16.785 ;
        RECT 32.485 16.615 32.655 16.785 ;
        RECT 32.945 16.615 33.115 16.785 ;
        RECT 33.405 16.615 33.575 16.785 ;
        RECT 33.865 16.615 34.035 16.785 ;
        RECT 34.325 16.615 34.495 16.785 ;
        RECT 34.785 16.615 34.955 16.785 ;
        RECT 35.245 16.615 35.415 16.785 ;
        RECT 35.705 16.615 35.875 16.785 ;
        RECT 36.165 16.615 36.335 16.785 ;
        RECT 36.625 16.615 36.795 16.785 ;
        RECT 37.085 16.615 37.255 16.785 ;
        RECT 37.545 16.615 37.715 16.785 ;
        RECT 38.005 16.615 38.175 16.785 ;
        RECT 38.465 16.615 38.635 16.785 ;
        RECT 38.925 16.615 39.095 16.785 ;
        RECT 39.385 16.615 39.555 16.785 ;
        RECT 39.845 16.615 40.015 16.785 ;
        RECT 40.305 16.615 40.475 16.785 ;
        RECT 40.765 16.615 40.935 16.785 ;
        RECT 41.225 16.615 41.395 16.785 ;
        RECT 41.685 16.615 41.855 16.785 ;
        RECT 42.145 16.615 42.315 16.785 ;
        RECT 42.605 16.615 42.775 16.785 ;
        RECT 43.065 16.615 43.235 16.785 ;
        RECT 43.525 16.615 43.695 16.785 ;
        RECT 43.985 16.615 44.155 16.785 ;
        RECT 44.445 16.615 44.615 16.785 ;
        RECT 44.905 16.615 45.075 16.785 ;
        RECT 45.365 16.615 45.535 16.785 ;
        RECT 45.825 16.615 45.995 16.785 ;
        RECT 46.285 16.615 46.455 16.785 ;
        RECT 46.745 16.615 46.915 16.785 ;
        RECT 47.205 16.615 47.375 16.785 ;
        RECT 47.665 16.615 47.835 16.785 ;
        RECT 48.125 16.615 48.295 16.785 ;
        RECT 48.585 16.615 48.755 16.785 ;
        RECT 49.045 16.615 49.215 16.785 ;
        RECT 49.505 16.615 49.675 16.785 ;
        RECT 49.965 16.615 50.135 16.785 ;
        RECT 50.425 16.615 50.595 16.785 ;
        RECT 50.885 16.615 51.055 16.785 ;
        RECT 51.345 16.615 51.515 16.785 ;
        RECT 51.805 16.615 51.975 16.785 ;
        RECT 52.265 16.615 52.435 16.785 ;
        RECT 52.725 16.615 52.895 16.785 ;
        RECT 53.185 16.615 53.355 16.785 ;
        RECT 53.645 16.615 53.815 16.785 ;
        RECT 54.105 16.615 54.275 16.785 ;
        RECT 54.565 16.615 54.735 16.785 ;
        RECT 55.025 16.615 55.195 16.785 ;
        RECT 55.485 16.615 55.655 16.785 ;
        RECT 55.945 16.615 56.115 16.785 ;
        RECT 56.405 16.615 56.575 16.785 ;
        RECT 56.865 16.615 57.035 16.785 ;
        RECT 57.325 16.615 57.495 16.785 ;
        RECT 57.785 16.615 57.955 16.785 ;
        RECT 58.245 16.615 58.415 16.785 ;
        RECT 58.705 16.615 58.875 16.785 ;
        RECT 59.165 16.615 59.335 16.785 ;
        RECT 59.625 16.615 59.795 16.785 ;
        RECT 60.085 16.615 60.255 16.785 ;
        RECT 60.545 16.615 60.715 16.785 ;
        RECT 61.005 16.615 61.175 16.785 ;
        RECT 61.465 16.615 61.635 16.785 ;
        RECT 61.925 16.615 62.095 16.785 ;
        RECT 62.385 16.615 62.555 16.785 ;
        RECT 62.845 16.615 63.015 16.785 ;
        RECT 63.305 16.615 63.475 16.785 ;
        RECT 63.765 16.615 63.935 16.785 ;
        RECT 64.225 16.615 64.395 16.785 ;
        RECT 64.685 16.615 64.855 16.785 ;
        RECT 65.145 16.615 65.315 16.785 ;
        RECT 65.605 16.615 65.775 16.785 ;
        RECT 66.065 16.615 66.235 16.785 ;
        RECT 66.525 16.615 66.695 16.785 ;
        RECT 66.985 16.615 67.155 16.785 ;
        RECT 67.445 16.615 67.615 16.785 ;
        RECT 67.905 16.615 68.075 16.785 ;
        RECT 68.365 16.615 68.535 16.785 ;
        RECT 68.825 16.615 68.995 16.785 ;
        RECT 69.285 16.615 69.455 16.785 ;
        RECT 69.745 16.615 69.915 16.785 ;
        RECT 70.205 16.615 70.375 16.785 ;
        RECT 70.665 16.615 70.835 16.785 ;
        RECT 71.125 16.615 71.295 16.785 ;
        RECT 71.585 16.615 71.755 16.785 ;
        RECT 72.045 16.615 72.215 16.785 ;
        RECT 72.505 16.615 72.675 16.785 ;
        RECT 72.965 16.615 73.135 16.785 ;
        RECT 73.425 16.615 73.595 16.785 ;
        RECT 73.885 16.615 74.055 16.785 ;
        RECT 74.345 16.615 74.515 16.785 ;
        RECT 74.805 16.615 74.975 16.785 ;
        RECT 75.265 16.615 75.435 16.785 ;
        RECT 75.725 16.615 75.895 16.785 ;
        RECT 76.185 16.615 76.355 16.785 ;
        RECT 76.645 16.615 76.815 16.785 ;
        RECT 77.105 16.615 77.275 16.785 ;
        RECT 77.565 16.615 77.735 16.785 ;
        RECT 78.025 16.615 78.195 16.785 ;
        RECT 78.485 16.615 78.655 16.785 ;
        RECT 78.945 16.615 79.115 16.785 ;
        RECT 79.405 16.615 79.575 16.785 ;
        RECT 79.865 16.615 80.035 16.785 ;
        RECT 80.325 16.615 80.495 16.785 ;
        RECT 80.785 16.615 80.955 16.785 ;
        RECT 81.245 16.615 81.415 16.785 ;
        RECT 81.705 16.615 81.875 16.785 ;
        RECT 82.165 16.615 82.335 16.785 ;
        RECT 82.625 16.615 82.795 16.785 ;
        RECT 83.085 16.615 83.255 16.785 ;
        RECT 83.545 16.615 83.715 16.785 ;
        RECT 84.005 16.615 84.175 16.785 ;
        RECT 84.465 16.615 84.635 16.785 ;
        RECT 84.925 16.615 85.095 16.785 ;
        RECT 85.385 16.615 85.555 16.785 ;
        RECT 85.845 16.615 86.015 16.785 ;
        RECT 86.305 16.615 86.475 16.785 ;
        RECT 86.765 16.615 86.935 16.785 ;
        RECT 87.225 16.615 87.395 16.785 ;
        RECT 87.685 16.615 87.855 16.785 ;
        RECT 88.145 16.615 88.315 16.785 ;
        RECT 88.605 16.615 88.775 16.785 ;
        RECT 89.065 16.615 89.235 16.785 ;
        RECT 89.525 16.615 89.695 16.785 ;
        RECT 89.985 16.615 90.155 16.785 ;
        RECT 90.445 16.615 90.615 16.785 ;
        RECT 90.905 16.615 91.075 16.785 ;
        RECT 91.365 16.615 91.535 16.785 ;
        RECT 91.825 16.615 91.995 16.785 ;
        RECT 92.285 16.615 92.455 16.785 ;
        RECT 92.745 16.615 92.915 16.785 ;
        RECT 93.205 16.615 93.375 16.785 ;
        RECT 93.665 16.615 93.835 16.785 ;
        RECT 94.125 16.615 94.295 16.785 ;
        RECT 94.585 16.615 94.755 16.785 ;
        RECT 95.045 16.615 95.215 16.785 ;
        RECT 95.505 16.615 95.675 16.785 ;
        RECT 95.965 16.615 96.135 16.785 ;
        RECT 96.425 16.615 96.595 16.785 ;
        RECT 96.885 16.615 97.055 16.785 ;
        RECT 97.345 16.615 97.515 16.785 ;
        RECT 97.805 16.615 97.975 16.785 ;
        RECT 98.265 16.615 98.435 16.785 ;
        RECT 98.725 16.615 98.895 16.785 ;
        RECT 99.185 16.615 99.355 16.785 ;
        RECT 99.645 16.615 99.815 16.785 ;
      LAYER met1 ;
        RECT 16.700 98.060 99.960 98.540 ;
        RECT 16.700 92.620 99.960 93.100 ;
        RECT 16.700 87.180 99.960 87.660 ;
        RECT 16.700 81.740 99.960 82.220 ;
        RECT 16.700 76.300 99.960 76.780 ;
        RECT 16.700 70.860 99.960 71.340 ;
        RECT 16.700 65.420 99.960 65.900 ;
        RECT 16.700 59.980 99.960 60.460 ;
        RECT 16.700 54.540 99.960 55.020 ;
        RECT 16.700 49.100 99.960 49.580 ;
        RECT 16.700 43.660 99.960 44.140 ;
        RECT 16.700 38.220 99.960 38.700 ;
        RECT 16.700 32.780 99.960 33.260 ;
        RECT 16.700 27.340 99.960 27.820 ;
        RECT 16.700 21.900 99.960 22.380 ;
        RECT 16.700 16.460 99.960 16.940 ;
      LAYER via ;
        RECT 29.965 98.170 30.225 98.430 ;
        RECT 30.285 98.170 30.545 98.430 ;
        RECT 30.605 98.170 30.865 98.430 ;
        RECT 30.925 98.170 31.185 98.430 ;
        RECT 57.720 98.170 57.980 98.430 ;
        RECT 58.040 98.170 58.300 98.430 ;
        RECT 58.360 98.170 58.620 98.430 ;
        RECT 58.680 98.170 58.940 98.430 ;
        RECT 85.470 98.170 85.730 98.430 ;
        RECT 85.790 98.170 86.050 98.430 ;
        RECT 86.110 98.170 86.370 98.430 ;
        RECT 86.430 98.170 86.690 98.430 ;
        RECT 29.965 92.730 30.225 92.990 ;
        RECT 30.285 92.730 30.545 92.990 ;
        RECT 30.605 92.730 30.865 92.990 ;
        RECT 30.925 92.730 31.185 92.990 ;
        RECT 57.720 92.730 57.980 92.990 ;
        RECT 58.040 92.730 58.300 92.990 ;
        RECT 58.360 92.730 58.620 92.990 ;
        RECT 58.680 92.730 58.940 92.990 ;
        RECT 85.470 92.730 85.730 92.990 ;
        RECT 85.790 92.730 86.050 92.990 ;
        RECT 86.110 92.730 86.370 92.990 ;
        RECT 86.430 92.730 86.690 92.990 ;
        RECT 29.965 87.290 30.225 87.550 ;
        RECT 30.285 87.290 30.545 87.550 ;
        RECT 30.605 87.290 30.865 87.550 ;
        RECT 30.925 87.290 31.185 87.550 ;
        RECT 57.720 87.290 57.980 87.550 ;
        RECT 58.040 87.290 58.300 87.550 ;
        RECT 58.360 87.290 58.620 87.550 ;
        RECT 58.680 87.290 58.940 87.550 ;
        RECT 85.470 87.290 85.730 87.550 ;
        RECT 85.790 87.290 86.050 87.550 ;
        RECT 86.110 87.290 86.370 87.550 ;
        RECT 86.430 87.290 86.690 87.550 ;
        RECT 29.965 81.850 30.225 82.110 ;
        RECT 30.285 81.850 30.545 82.110 ;
        RECT 30.605 81.850 30.865 82.110 ;
        RECT 30.925 81.850 31.185 82.110 ;
        RECT 57.720 81.850 57.980 82.110 ;
        RECT 58.040 81.850 58.300 82.110 ;
        RECT 58.360 81.850 58.620 82.110 ;
        RECT 58.680 81.850 58.940 82.110 ;
        RECT 85.470 81.850 85.730 82.110 ;
        RECT 85.790 81.850 86.050 82.110 ;
        RECT 86.110 81.850 86.370 82.110 ;
        RECT 86.430 81.850 86.690 82.110 ;
        RECT 29.965 76.410 30.225 76.670 ;
        RECT 30.285 76.410 30.545 76.670 ;
        RECT 30.605 76.410 30.865 76.670 ;
        RECT 30.925 76.410 31.185 76.670 ;
        RECT 57.720 76.410 57.980 76.670 ;
        RECT 58.040 76.410 58.300 76.670 ;
        RECT 58.360 76.410 58.620 76.670 ;
        RECT 58.680 76.410 58.940 76.670 ;
        RECT 85.470 76.410 85.730 76.670 ;
        RECT 85.790 76.410 86.050 76.670 ;
        RECT 86.110 76.410 86.370 76.670 ;
        RECT 86.430 76.410 86.690 76.670 ;
        RECT 29.965 70.970 30.225 71.230 ;
        RECT 30.285 70.970 30.545 71.230 ;
        RECT 30.605 70.970 30.865 71.230 ;
        RECT 30.925 70.970 31.185 71.230 ;
        RECT 57.720 70.970 57.980 71.230 ;
        RECT 58.040 70.970 58.300 71.230 ;
        RECT 58.360 70.970 58.620 71.230 ;
        RECT 58.680 70.970 58.940 71.230 ;
        RECT 85.470 70.970 85.730 71.230 ;
        RECT 85.790 70.970 86.050 71.230 ;
        RECT 86.110 70.970 86.370 71.230 ;
        RECT 86.430 70.970 86.690 71.230 ;
        RECT 29.965 65.530 30.225 65.790 ;
        RECT 30.285 65.530 30.545 65.790 ;
        RECT 30.605 65.530 30.865 65.790 ;
        RECT 30.925 65.530 31.185 65.790 ;
        RECT 57.720 65.530 57.980 65.790 ;
        RECT 58.040 65.530 58.300 65.790 ;
        RECT 58.360 65.530 58.620 65.790 ;
        RECT 58.680 65.530 58.940 65.790 ;
        RECT 85.470 65.530 85.730 65.790 ;
        RECT 85.790 65.530 86.050 65.790 ;
        RECT 86.110 65.530 86.370 65.790 ;
        RECT 86.430 65.530 86.690 65.790 ;
        RECT 29.965 60.090 30.225 60.350 ;
        RECT 30.285 60.090 30.545 60.350 ;
        RECT 30.605 60.090 30.865 60.350 ;
        RECT 30.925 60.090 31.185 60.350 ;
        RECT 57.720 60.090 57.980 60.350 ;
        RECT 58.040 60.090 58.300 60.350 ;
        RECT 58.360 60.090 58.620 60.350 ;
        RECT 58.680 60.090 58.940 60.350 ;
        RECT 85.470 60.090 85.730 60.350 ;
        RECT 85.790 60.090 86.050 60.350 ;
        RECT 86.110 60.090 86.370 60.350 ;
        RECT 86.430 60.090 86.690 60.350 ;
        RECT 29.965 54.650 30.225 54.910 ;
        RECT 30.285 54.650 30.545 54.910 ;
        RECT 30.605 54.650 30.865 54.910 ;
        RECT 30.925 54.650 31.185 54.910 ;
        RECT 57.720 54.650 57.980 54.910 ;
        RECT 58.040 54.650 58.300 54.910 ;
        RECT 58.360 54.650 58.620 54.910 ;
        RECT 58.680 54.650 58.940 54.910 ;
        RECT 85.470 54.650 85.730 54.910 ;
        RECT 85.790 54.650 86.050 54.910 ;
        RECT 86.110 54.650 86.370 54.910 ;
        RECT 86.430 54.650 86.690 54.910 ;
        RECT 29.965 49.210 30.225 49.470 ;
        RECT 30.285 49.210 30.545 49.470 ;
        RECT 30.605 49.210 30.865 49.470 ;
        RECT 30.925 49.210 31.185 49.470 ;
        RECT 57.720 49.210 57.980 49.470 ;
        RECT 58.040 49.210 58.300 49.470 ;
        RECT 58.360 49.210 58.620 49.470 ;
        RECT 58.680 49.210 58.940 49.470 ;
        RECT 85.470 49.210 85.730 49.470 ;
        RECT 85.790 49.210 86.050 49.470 ;
        RECT 86.110 49.210 86.370 49.470 ;
        RECT 86.430 49.210 86.690 49.470 ;
        RECT 29.965 43.770 30.225 44.030 ;
        RECT 30.285 43.770 30.545 44.030 ;
        RECT 30.605 43.770 30.865 44.030 ;
        RECT 30.925 43.770 31.185 44.030 ;
        RECT 57.720 43.770 57.980 44.030 ;
        RECT 58.040 43.770 58.300 44.030 ;
        RECT 58.360 43.770 58.620 44.030 ;
        RECT 58.680 43.770 58.940 44.030 ;
        RECT 85.470 43.770 85.730 44.030 ;
        RECT 85.790 43.770 86.050 44.030 ;
        RECT 86.110 43.770 86.370 44.030 ;
        RECT 86.430 43.770 86.690 44.030 ;
        RECT 29.965 38.330 30.225 38.590 ;
        RECT 30.285 38.330 30.545 38.590 ;
        RECT 30.605 38.330 30.865 38.590 ;
        RECT 30.925 38.330 31.185 38.590 ;
        RECT 57.720 38.330 57.980 38.590 ;
        RECT 58.040 38.330 58.300 38.590 ;
        RECT 58.360 38.330 58.620 38.590 ;
        RECT 58.680 38.330 58.940 38.590 ;
        RECT 85.470 38.330 85.730 38.590 ;
        RECT 85.790 38.330 86.050 38.590 ;
        RECT 86.110 38.330 86.370 38.590 ;
        RECT 86.430 38.330 86.690 38.590 ;
        RECT 29.965 32.890 30.225 33.150 ;
        RECT 30.285 32.890 30.545 33.150 ;
        RECT 30.605 32.890 30.865 33.150 ;
        RECT 30.925 32.890 31.185 33.150 ;
        RECT 57.720 32.890 57.980 33.150 ;
        RECT 58.040 32.890 58.300 33.150 ;
        RECT 58.360 32.890 58.620 33.150 ;
        RECT 58.680 32.890 58.940 33.150 ;
        RECT 85.470 32.890 85.730 33.150 ;
        RECT 85.790 32.890 86.050 33.150 ;
        RECT 86.110 32.890 86.370 33.150 ;
        RECT 86.430 32.890 86.690 33.150 ;
        RECT 29.965 27.450 30.225 27.710 ;
        RECT 30.285 27.450 30.545 27.710 ;
        RECT 30.605 27.450 30.865 27.710 ;
        RECT 30.925 27.450 31.185 27.710 ;
        RECT 57.720 27.450 57.980 27.710 ;
        RECT 58.040 27.450 58.300 27.710 ;
        RECT 58.360 27.450 58.620 27.710 ;
        RECT 58.680 27.450 58.940 27.710 ;
        RECT 85.470 27.450 85.730 27.710 ;
        RECT 85.790 27.450 86.050 27.710 ;
        RECT 86.110 27.450 86.370 27.710 ;
        RECT 86.430 27.450 86.690 27.710 ;
        RECT 29.965 22.010 30.225 22.270 ;
        RECT 30.285 22.010 30.545 22.270 ;
        RECT 30.605 22.010 30.865 22.270 ;
        RECT 30.925 22.010 31.185 22.270 ;
        RECT 57.720 22.010 57.980 22.270 ;
        RECT 58.040 22.010 58.300 22.270 ;
        RECT 58.360 22.010 58.620 22.270 ;
        RECT 58.680 22.010 58.940 22.270 ;
        RECT 85.470 22.010 85.730 22.270 ;
        RECT 85.790 22.010 86.050 22.270 ;
        RECT 86.110 22.010 86.370 22.270 ;
        RECT 86.430 22.010 86.690 22.270 ;
        RECT 29.965 16.570 30.225 16.830 ;
        RECT 30.285 16.570 30.545 16.830 ;
        RECT 30.605 16.570 30.865 16.830 ;
        RECT 30.925 16.570 31.185 16.830 ;
        RECT 57.720 16.570 57.980 16.830 ;
        RECT 58.040 16.570 58.300 16.830 ;
        RECT 58.360 16.570 58.620 16.830 ;
        RECT 58.680 16.570 58.940 16.830 ;
        RECT 85.470 16.570 85.730 16.830 ;
        RECT 85.790 16.570 86.050 16.830 ;
        RECT 86.110 16.570 86.370 16.830 ;
        RECT 86.430 16.570 86.690 16.830 ;
      LAYER met2 ;
        RECT 29.835 98.060 31.315 98.540 ;
        RECT 57.590 98.060 59.070 98.540 ;
        RECT 85.340 98.060 86.820 98.540 ;
        RECT 29.835 92.620 31.315 93.100 ;
        RECT 57.590 92.620 59.070 93.100 ;
        RECT 85.340 92.620 86.820 93.100 ;
        RECT 29.835 87.180 31.315 87.660 ;
        RECT 57.590 87.180 59.070 87.660 ;
        RECT 85.340 87.180 86.820 87.660 ;
        RECT 29.835 81.740 31.315 82.220 ;
        RECT 57.590 81.740 59.070 82.220 ;
        RECT 85.340 81.740 86.820 82.220 ;
        RECT 29.835 76.300 31.315 76.780 ;
        RECT 57.590 76.300 59.070 76.780 ;
        RECT 85.340 76.300 86.820 76.780 ;
        RECT 29.835 70.860 31.315 71.340 ;
        RECT 57.590 70.860 59.070 71.340 ;
        RECT 85.340 70.860 86.820 71.340 ;
        RECT 29.835 65.420 31.315 65.900 ;
        RECT 57.590 65.420 59.070 65.900 ;
        RECT 85.340 65.420 86.820 65.900 ;
        RECT 29.835 59.980 31.315 60.460 ;
        RECT 57.590 59.980 59.070 60.460 ;
        RECT 85.340 59.980 86.820 60.460 ;
        RECT 29.835 54.540 31.315 55.020 ;
        RECT 57.590 54.540 59.070 55.020 ;
        RECT 85.340 54.540 86.820 55.020 ;
        RECT 29.835 49.100 31.315 49.580 ;
        RECT 57.590 49.100 59.070 49.580 ;
        RECT 85.340 49.100 86.820 49.580 ;
        RECT 29.835 43.660 31.315 44.140 ;
        RECT 57.590 43.660 59.070 44.140 ;
        RECT 85.340 43.660 86.820 44.140 ;
        RECT 29.835 38.220 31.315 38.700 ;
        RECT 57.590 38.220 59.070 38.700 ;
        RECT 85.340 38.220 86.820 38.700 ;
        RECT 29.835 32.780 31.315 33.260 ;
        RECT 57.590 32.780 59.070 33.260 ;
        RECT 85.340 32.780 86.820 33.260 ;
        RECT 29.835 27.340 31.315 27.820 ;
        RECT 57.590 27.340 59.070 27.820 ;
        RECT 85.340 27.340 86.820 27.820 ;
        RECT 29.835 21.900 31.315 22.380 ;
        RECT 57.590 21.900 59.070 22.380 ;
        RECT 85.340 21.900 86.820 22.380 ;
        RECT 29.835 16.460 31.315 16.940 ;
        RECT 57.590 16.460 59.070 16.940 ;
        RECT 85.340 16.460 86.820 16.940 ;
      LAYER via2 ;
        RECT 29.835 98.160 30.115 98.440 ;
        RECT 30.235 98.160 30.515 98.440 ;
        RECT 30.635 98.160 30.915 98.440 ;
        RECT 31.035 98.160 31.315 98.440 ;
        RECT 57.590 98.160 57.870 98.440 ;
        RECT 57.990 98.160 58.270 98.440 ;
        RECT 58.390 98.160 58.670 98.440 ;
        RECT 58.790 98.160 59.070 98.440 ;
        RECT 85.340 98.160 85.620 98.440 ;
        RECT 85.740 98.160 86.020 98.440 ;
        RECT 86.140 98.160 86.420 98.440 ;
        RECT 86.540 98.160 86.820 98.440 ;
        RECT 29.835 92.720 30.115 93.000 ;
        RECT 30.235 92.720 30.515 93.000 ;
        RECT 30.635 92.720 30.915 93.000 ;
        RECT 31.035 92.720 31.315 93.000 ;
        RECT 57.590 92.720 57.870 93.000 ;
        RECT 57.990 92.720 58.270 93.000 ;
        RECT 58.390 92.720 58.670 93.000 ;
        RECT 58.790 92.720 59.070 93.000 ;
        RECT 85.340 92.720 85.620 93.000 ;
        RECT 85.740 92.720 86.020 93.000 ;
        RECT 86.140 92.720 86.420 93.000 ;
        RECT 86.540 92.720 86.820 93.000 ;
        RECT 29.835 87.280 30.115 87.560 ;
        RECT 30.235 87.280 30.515 87.560 ;
        RECT 30.635 87.280 30.915 87.560 ;
        RECT 31.035 87.280 31.315 87.560 ;
        RECT 57.590 87.280 57.870 87.560 ;
        RECT 57.990 87.280 58.270 87.560 ;
        RECT 58.390 87.280 58.670 87.560 ;
        RECT 58.790 87.280 59.070 87.560 ;
        RECT 85.340 87.280 85.620 87.560 ;
        RECT 85.740 87.280 86.020 87.560 ;
        RECT 86.140 87.280 86.420 87.560 ;
        RECT 86.540 87.280 86.820 87.560 ;
        RECT 29.835 81.840 30.115 82.120 ;
        RECT 30.235 81.840 30.515 82.120 ;
        RECT 30.635 81.840 30.915 82.120 ;
        RECT 31.035 81.840 31.315 82.120 ;
        RECT 57.590 81.840 57.870 82.120 ;
        RECT 57.990 81.840 58.270 82.120 ;
        RECT 58.390 81.840 58.670 82.120 ;
        RECT 58.790 81.840 59.070 82.120 ;
        RECT 85.340 81.840 85.620 82.120 ;
        RECT 85.740 81.840 86.020 82.120 ;
        RECT 86.140 81.840 86.420 82.120 ;
        RECT 86.540 81.840 86.820 82.120 ;
        RECT 29.835 76.400 30.115 76.680 ;
        RECT 30.235 76.400 30.515 76.680 ;
        RECT 30.635 76.400 30.915 76.680 ;
        RECT 31.035 76.400 31.315 76.680 ;
        RECT 57.590 76.400 57.870 76.680 ;
        RECT 57.990 76.400 58.270 76.680 ;
        RECT 58.390 76.400 58.670 76.680 ;
        RECT 58.790 76.400 59.070 76.680 ;
        RECT 85.340 76.400 85.620 76.680 ;
        RECT 85.740 76.400 86.020 76.680 ;
        RECT 86.140 76.400 86.420 76.680 ;
        RECT 86.540 76.400 86.820 76.680 ;
        RECT 29.835 70.960 30.115 71.240 ;
        RECT 30.235 70.960 30.515 71.240 ;
        RECT 30.635 70.960 30.915 71.240 ;
        RECT 31.035 70.960 31.315 71.240 ;
        RECT 57.590 70.960 57.870 71.240 ;
        RECT 57.990 70.960 58.270 71.240 ;
        RECT 58.390 70.960 58.670 71.240 ;
        RECT 58.790 70.960 59.070 71.240 ;
        RECT 85.340 70.960 85.620 71.240 ;
        RECT 85.740 70.960 86.020 71.240 ;
        RECT 86.140 70.960 86.420 71.240 ;
        RECT 86.540 70.960 86.820 71.240 ;
        RECT 29.835 65.520 30.115 65.800 ;
        RECT 30.235 65.520 30.515 65.800 ;
        RECT 30.635 65.520 30.915 65.800 ;
        RECT 31.035 65.520 31.315 65.800 ;
        RECT 57.590 65.520 57.870 65.800 ;
        RECT 57.990 65.520 58.270 65.800 ;
        RECT 58.390 65.520 58.670 65.800 ;
        RECT 58.790 65.520 59.070 65.800 ;
        RECT 85.340 65.520 85.620 65.800 ;
        RECT 85.740 65.520 86.020 65.800 ;
        RECT 86.140 65.520 86.420 65.800 ;
        RECT 86.540 65.520 86.820 65.800 ;
        RECT 29.835 60.080 30.115 60.360 ;
        RECT 30.235 60.080 30.515 60.360 ;
        RECT 30.635 60.080 30.915 60.360 ;
        RECT 31.035 60.080 31.315 60.360 ;
        RECT 57.590 60.080 57.870 60.360 ;
        RECT 57.990 60.080 58.270 60.360 ;
        RECT 58.390 60.080 58.670 60.360 ;
        RECT 58.790 60.080 59.070 60.360 ;
        RECT 85.340 60.080 85.620 60.360 ;
        RECT 85.740 60.080 86.020 60.360 ;
        RECT 86.140 60.080 86.420 60.360 ;
        RECT 86.540 60.080 86.820 60.360 ;
        RECT 29.835 54.640 30.115 54.920 ;
        RECT 30.235 54.640 30.515 54.920 ;
        RECT 30.635 54.640 30.915 54.920 ;
        RECT 31.035 54.640 31.315 54.920 ;
        RECT 57.590 54.640 57.870 54.920 ;
        RECT 57.990 54.640 58.270 54.920 ;
        RECT 58.390 54.640 58.670 54.920 ;
        RECT 58.790 54.640 59.070 54.920 ;
        RECT 85.340 54.640 85.620 54.920 ;
        RECT 85.740 54.640 86.020 54.920 ;
        RECT 86.140 54.640 86.420 54.920 ;
        RECT 86.540 54.640 86.820 54.920 ;
        RECT 29.835 49.200 30.115 49.480 ;
        RECT 30.235 49.200 30.515 49.480 ;
        RECT 30.635 49.200 30.915 49.480 ;
        RECT 31.035 49.200 31.315 49.480 ;
        RECT 57.590 49.200 57.870 49.480 ;
        RECT 57.990 49.200 58.270 49.480 ;
        RECT 58.390 49.200 58.670 49.480 ;
        RECT 58.790 49.200 59.070 49.480 ;
        RECT 85.340 49.200 85.620 49.480 ;
        RECT 85.740 49.200 86.020 49.480 ;
        RECT 86.140 49.200 86.420 49.480 ;
        RECT 86.540 49.200 86.820 49.480 ;
        RECT 29.835 43.760 30.115 44.040 ;
        RECT 30.235 43.760 30.515 44.040 ;
        RECT 30.635 43.760 30.915 44.040 ;
        RECT 31.035 43.760 31.315 44.040 ;
        RECT 57.590 43.760 57.870 44.040 ;
        RECT 57.990 43.760 58.270 44.040 ;
        RECT 58.390 43.760 58.670 44.040 ;
        RECT 58.790 43.760 59.070 44.040 ;
        RECT 85.340 43.760 85.620 44.040 ;
        RECT 85.740 43.760 86.020 44.040 ;
        RECT 86.140 43.760 86.420 44.040 ;
        RECT 86.540 43.760 86.820 44.040 ;
        RECT 29.835 38.320 30.115 38.600 ;
        RECT 30.235 38.320 30.515 38.600 ;
        RECT 30.635 38.320 30.915 38.600 ;
        RECT 31.035 38.320 31.315 38.600 ;
        RECT 57.590 38.320 57.870 38.600 ;
        RECT 57.990 38.320 58.270 38.600 ;
        RECT 58.390 38.320 58.670 38.600 ;
        RECT 58.790 38.320 59.070 38.600 ;
        RECT 85.340 38.320 85.620 38.600 ;
        RECT 85.740 38.320 86.020 38.600 ;
        RECT 86.140 38.320 86.420 38.600 ;
        RECT 86.540 38.320 86.820 38.600 ;
        RECT 29.835 32.880 30.115 33.160 ;
        RECT 30.235 32.880 30.515 33.160 ;
        RECT 30.635 32.880 30.915 33.160 ;
        RECT 31.035 32.880 31.315 33.160 ;
        RECT 57.590 32.880 57.870 33.160 ;
        RECT 57.990 32.880 58.270 33.160 ;
        RECT 58.390 32.880 58.670 33.160 ;
        RECT 58.790 32.880 59.070 33.160 ;
        RECT 85.340 32.880 85.620 33.160 ;
        RECT 85.740 32.880 86.020 33.160 ;
        RECT 86.140 32.880 86.420 33.160 ;
        RECT 86.540 32.880 86.820 33.160 ;
        RECT 29.835 27.440 30.115 27.720 ;
        RECT 30.235 27.440 30.515 27.720 ;
        RECT 30.635 27.440 30.915 27.720 ;
        RECT 31.035 27.440 31.315 27.720 ;
        RECT 57.590 27.440 57.870 27.720 ;
        RECT 57.990 27.440 58.270 27.720 ;
        RECT 58.390 27.440 58.670 27.720 ;
        RECT 58.790 27.440 59.070 27.720 ;
        RECT 85.340 27.440 85.620 27.720 ;
        RECT 85.740 27.440 86.020 27.720 ;
        RECT 86.140 27.440 86.420 27.720 ;
        RECT 86.540 27.440 86.820 27.720 ;
        RECT 29.835 22.000 30.115 22.280 ;
        RECT 30.235 22.000 30.515 22.280 ;
        RECT 30.635 22.000 30.915 22.280 ;
        RECT 31.035 22.000 31.315 22.280 ;
        RECT 57.590 22.000 57.870 22.280 ;
        RECT 57.990 22.000 58.270 22.280 ;
        RECT 58.390 22.000 58.670 22.280 ;
        RECT 58.790 22.000 59.070 22.280 ;
        RECT 85.340 22.000 85.620 22.280 ;
        RECT 85.740 22.000 86.020 22.280 ;
        RECT 86.140 22.000 86.420 22.280 ;
        RECT 86.540 22.000 86.820 22.280 ;
        RECT 29.835 16.560 30.115 16.840 ;
        RECT 30.235 16.560 30.515 16.840 ;
        RECT 30.635 16.560 30.915 16.840 ;
        RECT 31.035 16.560 31.315 16.840 ;
        RECT 57.590 16.560 57.870 16.840 ;
        RECT 57.990 16.560 58.270 16.840 ;
        RECT 58.390 16.560 58.670 16.840 ;
        RECT 58.790 16.560 59.070 16.840 ;
        RECT 85.340 16.560 85.620 16.840 ;
        RECT 85.740 16.560 86.020 16.840 ;
        RECT 86.140 16.560 86.420 16.840 ;
        RECT 86.540 16.560 86.820 16.840 ;
      LAYER met3 ;
        RECT 29.775 98.135 31.375 98.465 ;
        RECT 57.530 98.135 59.130 98.465 ;
        RECT 85.280 98.135 86.880 98.465 ;
        RECT 29.775 92.695 31.375 93.025 ;
        RECT 57.530 92.695 59.130 93.025 ;
        RECT 85.280 92.695 86.880 93.025 ;
        RECT 29.775 87.255 31.375 87.585 ;
        RECT 57.530 87.255 59.130 87.585 ;
        RECT 85.280 87.255 86.880 87.585 ;
        RECT 29.775 81.815 31.375 82.145 ;
        RECT 57.530 81.815 59.130 82.145 ;
        RECT 85.280 81.815 86.880 82.145 ;
        RECT 29.775 76.375 31.375 76.705 ;
        RECT 57.530 76.375 59.130 76.705 ;
        RECT 85.280 76.375 86.880 76.705 ;
        RECT 29.775 70.935 31.375 71.265 ;
        RECT 57.530 70.935 59.130 71.265 ;
        RECT 85.280 70.935 86.880 71.265 ;
        RECT 29.775 65.495 31.375 65.825 ;
        RECT 57.530 65.495 59.130 65.825 ;
        RECT 85.280 65.495 86.880 65.825 ;
        RECT 29.775 60.055 31.375 60.385 ;
        RECT 57.530 60.055 59.130 60.385 ;
        RECT 85.280 60.055 86.880 60.385 ;
        RECT 29.775 54.615 31.375 54.945 ;
        RECT 57.530 54.615 59.130 54.945 ;
        RECT 85.280 54.615 86.880 54.945 ;
        RECT 29.775 49.175 31.375 49.505 ;
        RECT 57.530 49.175 59.130 49.505 ;
        RECT 85.280 49.175 86.880 49.505 ;
        RECT 29.775 43.735 31.375 44.065 ;
        RECT 57.530 43.735 59.130 44.065 ;
        RECT 85.280 43.735 86.880 44.065 ;
        RECT 29.775 38.295 31.375 38.625 ;
        RECT 57.530 38.295 59.130 38.625 ;
        RECT 85.280 38.295 86.880 38.625 ;
        RECT 29.775 32.855 31.375 33.185 ;
        RECT 57.530 32.855 59.130 33.185 ;
        RECT 85.280 32.855 86.880 33.185 ;
        RECT 29.775 27.415 31.375 27.745 ;
        RECT 57.530 27.415 59.130 27.745 ;
        RECT 85.280 27.415 86.880 27.745 ;
        RECT 29.775 21.975 31.375 22.305 ;
        RECT 57.530 21.975 59.130 22.305 ;
        RECT 85.280 21.975 86.880 22.305 ;
        RECT 29.775 16.535 31.375 16.865 ;
        RECT 57.530 16.535 59.130 16.865 ;
        RECT 85.280 16.535 86.880 16.865 ;
      LAYER via3 ;
        RECT 29.815 98.140 30.135 98.460 ;
        RECT 30.215 98.140 30.535 98.460 ;
        RECT 30.615 98.140 30.935 98.460 ;
        RECT 31.015 98.140 31.335 98.460 ;
        RECT 57.570 98.140 57.890 98.460 ;
        RECT 57.970 98.140 58.290 98.460 ;
        RECT 58.370 98.140 58.690 98.460 ;
        RECT 58.770 98.140 59.090 98.460 ;
        RECT 85.320 98.140 85.640 98.460 ;
        RECT 85.720 98.140 86.040 98.460 ;
        RECT 86.120 98.140 86.440 98.460 ;
        RECT 86.520 98.140 86.840 98.460 ;
        RECT 29.815 92.700 30.135 93.020 ;
        RECT 30.215 92.700 30.535 93.020 ;
        RECT 30.615 92.700 30.935 93.020 ;
        RECT 31.015 92.700 31.335 93.020 ;
        RECT 57.570 92.700 57.890 93.020 ;
        RECT 57.970 92.700 58.290 93.020 ;
        RECT 58.370 92.700 58.690 93.020 ;
        RECT 58.770 92.700 59.090 93.020 ;
        RECT 85.320 92.700 85.640 93.020 ;
        RECT 85.720 92.700 86.040 93.020 ;
        RECT 86.120 92.700 86.440 93.020 ;
        RECT 86.520 92.700 86.840 93.020 ;
        RECT 29.815 87.260 30.135 87.580 ;
        RECT 30.215 87.260 30.535 87.580 ;
        RECT 30.615 87.260 30.935 87.580 ;
        RECT 31.015 87.260 31.335 87.580 ;
        RECT 57.570 87.260 57.890 87.580 ;
        RECT 57.970 87.260 58.290 87.580 ;
        RECT 58.370 87.260 58.690 87.580 ;
        RECT 58.770 87.260 59.090 87.580 ;
        RECT 85.320 87.260 85.640 87.580 ;
        RECT 85.720 87.260 86.040 87.580 ;
        RECT 86.120 87.260 86.440 87.580 ;
        RECT 86.520 87.260 86.840 87.580 ;
        RECT 29.815 81.820 30.135 82.140 ;
        RECT 30.215 81.820 30.535 82.140 ;
        RECT 30.615 81.820 30.935 82.140 ;
        RECT 31.015 81.820 31.335 82.140 ;
        RECT 57.570 81.820 57.890 82.140 ;
        RECT 57.970 81.820 58.290 82.140 ;
        RECT 58.370 81.820 58.690 82.140 ;
        RECT 58.770 81.820 59.090 82.140 ;
        RECT 85.320 81.820 85.640 82.140 ;
        RECT 85.720 81.820 86.040 82.140 ;
        RECT 86.120 81.820 86.440 82.140 ;
        RECT 86.520 81.820 86.840 82.140 ;
        RECT 29.815 76.380 30.135 76.700 ;
        RECT 30.215 76.380 30.535 76.700 ;
        RECT 30.615 76.380 30.935 76.700 ;
        RECT 31.015 76.380 31.335 76.700 ;
        RECT 57.570 76.380 57.890 76.700 ;
        RECT 57.970 76.380 58.290 76.700 ;
        RECT 58.370 76.380 58.690 76.700 ;
        RECT 58.770 76.380 59.090 76.700 ;
        RECT 85.320 76.380 85.640 76.700 ;
        RECT 85.720 76.380 86.040 76.700 ;
        RECT 86.120 76.380 86.440 76.700 ;
        RECT 86.520 76.380 86.840 76.700 ;
        RECT 29.815 70.940 30.135 71.260 ;
        RECT 30.215 70.940 30.535 71.260 ;
        RECT 30.615 70.940 30.935 71.260 ;
        RECT 31.015 70.940 31.335 71.260 ;
        RECT 57.570 70.940 57.890 71.260 ;
        RECT 57.970 70.940 58.290 71.260 ;
        RECT 58.370 70.940 58.690 71.260 ;
        RECT 58.770 70.940 59.090 71.260 ;
        RECT 85.320 70.940 85.640 71.260 ;
        RECT 85.720 70.940 86.040 71.260 ;
        RECT 86.120 70.940 86.440 71.260 ;
        RECT 86.520 70.940 86.840 71.260 ;
        RECT 29.815 65.500 30.135 65.820 ;
        RECT 30.215 65.500 30.535 65.820 ;
        RECT 30.615 65.500 30.935 65.820 ;
        RECT 31.015 65.500 31.335 65.820 ;
        RECT 57.570 65.500 57.890 65.820 ;
        RECT 57.970 65.500 58.290 65.820 ;
        RECT 58.370 65.500 58.690 65.820 ;
        RECT 58.770 65.500 59.090 65.820 ;
        RECT 85.320 65.500 85.640 65.820 ;
        RECT 85.720 65.500 86.040 65.820 ;
        RECT 86.120 65.500 86.440 65.820 ;
        RECT 86.520 65.500 86.840 65.820 ;
        RECT 29.815 60.060 30.135 60.380 ;
        RECT 30.215 60.060 30.535 60.380 ;
        RECT 30.615 60.060 30.935 60.380 ;
        RECT 31.015 60.060 31.335 60.380 ;
        RECT 57.570 60.060 57.890 60.380 ;
        RECT 57.970 60.060 58.290 60.380 ;
        RECT 58.370 60.060 58.690 60.380 ;
        RECT 58.770 60.060 59.090 60.380 ;
        RECT 85.320 60.060 85.640 60.380 ;
        RECT 85.720 60.060 86.040 60.380 ;
        RECT 86.120 60.060 86.440 60.380 ;
        RECT 86.520 60.060 86.840 60.380 ;
        RECT 29.815 54.620 30.135 54.940 ;
        RECT 30.215 54.620 30.535 54.940 ;
        RECT 30.615 54.620 30.935 54.940 ;
        RECT 31.015 54.620 31.335 54.940 ;
        RECT 57.570 54.620 57.890 54.940 ;
        RECT 57.970 54.620 58.290 54.940 ;
        RECT 58.370 54.620 58.690 54.940 ;
        RECT 58.770 54.620 59.090 54.940 ;
        RECT 85.320 54.620 85.640 54.940 ;
        RECT 85.720 54.620 86.040 54.940 ;
        RECT 86.120 54.620 86.440 54.940 ;
        RECT 86.520 54.620 86.840 54.940 ;
        RECT 29.815 49.180 30.135 49.500 ;
        RECT 30.215 49.180 30.535 49.500 ;
        RECT 30.615 49.180 30.935 49.500 ;
        RECT 31.015 49.180 31.335 49.500 ;
        RECT 57.570 49.180 57.890 49.500 ;
        RECT 57.970 49.180 58.290 49.500 ;
        RECT 58.370 49.180 58.690 49.500 ;
        RECT 58.770 49.180 59.090 49.500 ;
        RECT 85.320 49.180 85.640 49.500 ;
        RECT 85.720 49.180 86.040 49.500 ;
        RECT 86.120 49.180 86.440 49.500 ;
        RECT 86.520 49.180 86.840 49.500 ;
        RECT 29.815 43.740 30.135 44.060 ;
        RECT 30.215 43.740 30.535 44.060 ;
        RECT 30.615 43.740 30.935 44.060 ;
        RECT 31.015 43.740 31.335 44.060 ;
        RECT 57.570 43.740 57.890 44.060 ;
        RECT 57.970 43.740 58.290 44.060 ;
        RECT 58.370 43.740 58.690 44.060 ;
        RECT 58.770 43.740 59.090 44.060 ;
        RECT 85.320 43.740 85.640 44.060 ;
        RECT 85.720 43.740 86.040 44.060 ;
        RECT 86.120 43.740 86.440 44.060 ;
        RECT 86.520 43.740 86.840 44.060 ;
        RECT 29.815 38.300 30.135 38.620 ;
        RECT 30.215 38.300 30.535 38.620 ;
        RECT 30.615 38.300 30.935 38.620 ;
        RECT 31.015 38.300 31.335 38.620 ;
        RECT 57.570 38.300 57.890 38.620 ;
        RECT 57.970 38.300 58.290 38.620 ;
        RECT 58.370 38.300 58.690 38.620 ;
        RECT 58.770 38.300 59.090 38.620 ;
        RECT 85.320 38.300 85.640 38.620 ;
        RECT 85.720 38.300 86.040 38.620 ;
        RECT 86.120 38.300 86.440 38.620 ;
        RECT 86.520 38.300 86.840 38.620 ;
        RECT 29.815 32.860 30.135 33.180 ;
        RECT 30.215 32.860 30.535 33.180 ;
        RECT 30.615 32.860 30.935 33.180 ;
        RECT 31.015 32.860 31.335 33.180 ;
        RECT 57.570 32.860 57.890 33.180 ;
        RECT 57.970 32.860 58.290 33.180 ;
        RECT 58.370 32.860 58.690 33.180 ;
        RECT 58.770 32.860 59.090 33.180 ;
        RECT 85.320 32.860 85.640 33.180 ;
        RECT 85.720 32.860 86.040 33.180 ;
        RECT 86.120 32.860 86.440 33.180 ;
        RECT 86.520 32.860 86.840 33.180 ;
        RECT 29.815 27.420 30.135 27.740 ;
        RECT 30.215 27.420 30.535 27.740 ;
        RECT 30.615 27.420 30.935 27.740 ;
        RECT 31.015 27.420 31.335 27.740 ;
        RECT 57.570 27.420 57.890 27.740 ;
        RECT 57.970 27.420 58.290 27.740 ;
        RECT 58.370 27.420 58.690 27.740 ;
        RECT 58.770 27.420 59.090 27.740 ;
        RECT 85.320 27.420 85.640 27.740 ;
        RECT 85.720 27.420 86.040 27.740 ;
        RECT 86.120 27.420 86.440 27.740 ;
        RECT 86.520 27.420 86.840 27.740 ;
        RECT 29.815 21.980 30.135 22.300 ;
        RECT 30.215 21.980 30.535 22.300 ;
        RECT 30.615 21.980 30.935 22.300 ;
        RECT 31.015 21.980 31.335 22.300 ;
        RECT 57.570 21.980 57.890 22.300 ;
        RECT 57.970 21.980 58.290 22.300 ;
        RECT 58.370 21.980 58.690 22.300 ;
        RECT 58.770 21.980 59.090 22.300 ;
        RECT 85.320 21.980 85.640 22.300 ;
        RECT 85.720 21.980 86.040 22.300 ;
        RECT 86.120 21.980 86.440 22.300 ;
        RECT 86.520 21.980 86.840 22.300 ;
        RECT 29.815 16.540 30.135 16.860 ;
        RECT 30.215 16.540 30.535 16.860 ;
        RECT 30.615 16.540 30.935 16.860 ;
        RECT 31.015 16.540 31.335 16.860 ;
        RECT 57.570 16.540 57.890 16.860 ;
        RECT 57.970 16.540 58.290 16.860 ;
        RECT 58.370 16.540 58.690 16.860 ;
        RECT 58.770 16.540 59.090 16.860 ;
        RECT 85.320 16.540 85.640 16.860 ;
        RECT 85.720 16.540 86.040 16.860 ;
        RECT 86.120 16.540 86.440 16.860 ;
        RECT 86.520 16.540 86.840 16.860 ;
      LAYER met4 ;
        RECT 9.900 9.900 11.500 105.100 ;
        RECT 29.775 6.600 31.375 108.400 ;
        RECT 57.530 6.600 59.130 108.400 ;
        RECT 85.280 6.600 86.885 108.400 ;
        RECT 105.160 9.900 106.760 105.100 ;
      LAYER via4 ;
        RECT 10.110 103.710 11.290 104.890 ;
        RECT 10.110 83.870 11.290 85.050 ;
        RECT 10.110 56.670 11.290 57.850 ;
        RECT 10.110 29.470 11.290 30.650 ;
        RECT 10.110 10.110 11.290 11.290 ;
        RECT 29.985 103.710 31.165 104.890 ;
        RECT 29.985 83.870 31.165 85.050 ;
        RECT 29.985 56.670 31.165 57.850 ;
        RECT 29.985 29.470 31.165 30.650 ;
        RECT 29.985 10.110 31.165 11.290 ;
        RECT 57.740 103.710 58.920 104.890 ;
        RECT 57.740 83.870 58.920 85.050 ;
        RECT 57.740 56.670 58.920 57.850 ;
        RECT 57.740 29.470 58.920 30.650 ;
        RECT 57.740 10.110 58.920 11.290 ;
        RECT 85.490 103.710 86.670 104.890 ;
        RECT 85.490 83.870 86.670 85.050 ;
        RECT 85.490 56.670 86.670 57.850 ;
        RECT 85.490 29.470 86.670 30.650 ;
        RECT 85.490 10.110 86.670 11.290 ;
        RECT 105.370 103.710 106.550 104.890 ;
        RECT 105.370 83.870 106.550 85.050 ;
        RECT 105.370 56.670 106.550 57.850 ;
        RECT 105.370 29.470 106.550 30.650 ;
        RECT 105.370 10.110 106.550 11.290 ;
      LAYER met5 ;
        RECT 9.900 103.500 106.760 105.100 ;
        RECT 6.600 83.660 110.060 85.260 ;
        RECT 6.600 56.460 110.060 58.060 ;
        RECT 6.600 29.260 110.060 30.860 ;
        RECT 9.900 9.900 106.760 11.500 ;
    END
  END vccd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 16.845 95.495 17.015 95.665 ;
        RECT 17.305 95.495 17.475 95.665 ;
        RECT 17.765 95.495 17.935 95.665 ;
        RECT 18.225 95.495 18.395 95.665 ;
        RECT 18.685 95.495 18.855 95.665 ;
        RECT 19.145 95.495 19.315 95.665 ;
        RECT 19.605 95.495 19.775 95.665 ;
        RECT 20.065 95.495 20.235 95.665 ;
        RECT 20.525 95.495 20.695 95.665 ;
        RECT 20.985 95.495 21.155 95.665 ;
        RECT 21.445 95.495 21.615 95.665 ;
        RECT 21.905 95.495 22.075 95.665 ;
        RECT 22.365 95.495 22.535 95.665 ;
        RECT 22.825 95.495 22.995 95.665 ;
        RECT 23.285 95.495 23.455 95.665 ;
        RECT 23.745 95.495 23.915 95.665 ;
        RECT 24.205 95.495 24.375 95.665 ;
        RECT 24.665 95.495 24.835 95.665 ;
        RECT 25.125 95.495 25.295 95.665 ;
        RECT 25.585 95.495 25.755 95.665 ;
        RECT 26.045 95.495 26.215 95.665 ;
        RECT 26.505 95.495 26.675 95.665 ;
        RECT 26.965 95.495 27.135 95.665 ;
        RECT 27.425 95.495 27.595 95.665 ;
        RECT 27.885 95.495 28.055 95.665 ;
        RECT 28.345 95.495 28.515 95.665 ;
        RECT 28.805 95.495 28.975 95.665 ;
        RECT 29.265 95.495 29.435 95.665 ;
        RECT 29.725 95.495 29.895 95.665 ;
        RECT 30.185 95.495 30.355 95.665 ;
        RECT 30.645 95.495 30.815 95.665 ;
        RECT 31.105 95.495 31.275 95.665 ;
        RECT 31.565 95.495 31.735 95.665 ;
        RECT 32.025 95.495 32.195 95.665 ;
        RECT 32.485 95.495 32.655 95.665 ;
        RECT 32.945 95.495 33.115 95.665 ;
        RECT 33.405 95.495 33.575 95.665 ;
        RECT 33.865 95.495 34.035 95.665 ;
        RECT 34.325 95.495 34.495 95.665 ;
        RECT 34.785 95.495 34.955 95.665 ;
        RECT 35.245 95.495 35.415 95.665 ;
        RECT 35.705 95.495 35.875 95.665 ;
        RECT 36.165 95.495 36.335 95.665 ;
        RECT 36.625 95.495 36.795 95.665 ;
        RECT 37.085 95.495 37.255 95.665 ;
        RECT 37.545 95.495 37.715 95.665 ;
        RECT 38.005 95.495 38.175 95.665 ;
        RECT 38.465 95.495 38.635 95.665 ;
        RECT 38.925 95.495 39.095 95.665 ;
        RECT 39.385 95.495 39.555 95.665 ;
        RECT 39.845 95.495 40.015 95.665 ;
        RECT 40.305 95.495 40.475 95.665 ;
        RECT 40.765 95.495 40.935 95.665 ;
        RECT 41.225 95.495 41.395 95.665 ;
        RECT 41.685 95.495 41.855 95.665 ;
        RECT 42.145 95.495 42.315 95.665 ;
        RECT 42.605 95.495 42.775 95.665 ;
        RECT 43.065 95.495 43.235 95.665 ;
        RECT 43.525 95.495 43.695 95.665 ;
        RECT 43.985 95.495 44.155 95.665 ;
        RECT 44.445 95.495 44.615 95.665 ;
        RECT 44.905 95.495 45.075 95.665 ;
        RECT 45.365 95.495 45.535 95.665 ;
        RECT 45.825 95.495 45.995 95.665 ;
        RECT 46.285 95.495 46.455 95.665 ;
        RECT 46.745 95.495 46.915 95.665 ;
        RECT 47.205 95.495 47.375 95.665 ;
        RECT 47.665 95.495 47.835 95.665 ;
        RECT 48.125 95.495 48.295 95.665 ;
        RECT 48.585 95.495 48.755 95.665 ;
        RECT 49.045 95.495 49.215 95.665 ;
        RECT 49.505 95.495 49.675 95.665 ;
        RECT 49.965 95.495 50.135 95.665 ;
        RECT 50.425 95.495 50.595 95.665 ;
        RECT 50.885 95.495 51.055 95.665 ;
        RECT 51.345 95.495 51.515 95.665 ;
        RECT 51.805 95.495 51.975 95.665 ;
        RECT 52.265 95.495 52.435 95.665 ;
        RECT 52.725 95.495 52.895 95.665 ;
        RECT 53.185 95.495 53.355 95.665 ;
        RECT 53.645 95.495 53.815 95.665 ;
        RECT 54.105 95.495 54.275 95.665 ;
        RECT 54.565 95.495 54.735 95.665 ;
        RECT 55.025 95.495 55.195 95.665 ;
        RECT 55.485 95.495 55.655 95.665 ;
        RECT 55.945 95.495 56.115 95.665 ;
        RECT 56.405 95.495 56.575 95.665 ;
        RECT 56.865 95.495 57.035 95.665 ;
        RECT 57.325 95.495 57.495 95.665 ;
        RECT 57.785 95.495 57.955 95.665 ;
        RECT 58.245 95.495 58.415 95.665 ;
        RECT 58.705 95.495 58.875 95.665 ;
        RECT 59.165 95.495 59.335 95.665 ;
        RECT 59.625 95.495 59.795 95.665 ;
        RECT 60.085 95.495 60.255 95.665 ;
        RECT 60.545 95.495 60.715 95.665 ;
        RECT 61.005 95.495 61.175 95.665 ;
        RECT 61.465 95.495 61.635 95.665 ;
        RECT 61.925 95.495 62.095 95.665 ;
        RECT 62.385 95.495 62.555 95.665 ;
        RECT 62.845 95.495 63.015 95.665 ;
        RECT 63.305 95.495 63.475 95.665 ;
        RECT 63.765 95.495 63.935 95.665 ;
        RECT 64.225 95.495 64.395 95.665 ;
        RECT 64.685 95.495 64.855 95.665 ;
        RECT 65.145 95.495 65.315 95.665 ;
        RECT 65.605 95.495 65.775 95.665 ;
        RECT 66.065 95.495 66.235 95.665 ;
        RECT 66.525 95.495 66.695 95.665 ;
        RECT 66.985 95.495 67.155 95.665 ;
        RECT 67.445 95.495 67.615 95.665 ;
        RECT 67.905 95.495 68.075 95.665 ;
        RECT 68.365 95.495 68.535 95.665 ;
        RECT 68.825 95.495 68.995 95.665 ;
        RECT 69.285 95.495 69.455 95.665 ;
        RECT 69.745 95.495 69.915 95.665 ;
        RECT 70.205 95.495 70.375 95.665 ;
        RECT 70.665 95.495 70.835 95.665 ;
        RECT 71.125 95.495 71.295 95.665 ;
        RECT 71.585 95.495 71.755 95.665 ;
        RECT 72.045 95.495 72.215 95.665 ;
        RECT 72.505 95.495 72.675 95.665 ;
        RECT 72.965 95.495 73.135 95.665 ;
        RECT 73.425 95.495 73.595 95.665 ;
        RECT 73.885 95.495 74.055 95.665 ;
        RECT 74.345 95.495 74.515 95.665 ;
        RECT 74.805 95.495 74.975 95.665 ;
        RECT 75.265 95.495 75.435 95.665 ;
        RECT 75.725 95.495 75.895 95.665 ;
        RECT 76.185 95.495 76.355 95.665 ;
        RECT 76.645 95.495 76.815 95.665 ;
        RECT 77.105 95.495 77.275 95.665 ;
        RECT 77.565 95.495 77.735 95.665 ;
        RECT 78.025 95.495 78.195 95.665 ;
        RECT 78.485 95.495 78.655 95.665 ;
        RECT 78.945 95.495 79.115 95.665 ;
        RECT 79.405 95.495 79.575 95.665 ;
        RECT 79.865 95.495 80.035 95.665 ;
        RECT 80.325 95.495 80.495 95.665 ;
        RECT 80.785 95.495 80.955 95.665 ;
        RECT 81.245 95.495 81.415 95.665 ;
        RECT 81.705 95.495 81.875 95.665 ;
        RECT 82.165 95.495 82.335 95.665 ;
        RECT 82.625 95.495 82.795 95.665 ;
        RECT 83.085 95.495 83.255 95.665 ;
        RECT 83.545 95.495 83.715 95.665 ;
        RECT 84.005 95.495 84.175 95.665 ;
        RECT 84.465 95.495 84.635 95.665 ;
        RECT 84.925 95.495 85.095 95.665 ;
        RECT 85.385 95.495 85.555 95.665 ;
        RECT 85.845 95.495 86.015 95.665 ;
        RECT 86.305 95.495 86.475 95.665 ;
        RECT 86.765 95.495 86.935 95.665 ;
        RECT 87.225 95.495 87.395 95.665 ;
        RECT 87.685 95.495 87.855 95.665 ;
        RECT 88.145 95.495 88.315 95.665 ;
        RECT 88.605 95.495 88.775 95.665 ;
        RECT 89.065 95.495 89.235 95.665 ;
        RECT 89.525 95.495 89.695 95.665 ;
        RECT 89.985 95.495 90.155 95.665 ;
        RECT 90.445 95.495 90.615 95.665 ;
        RECT 90.905 95.495 91.075 95.665 ;
        RECT 91.365 95.495 91.535 95.665 ;
        RECT 91.825 95.495 91.995 95.665 ;
        RECT 92.285 95.495 92.455 95.665 ;
        RECT 92.745 95.495 92.915 95.665 ;
        RECT 93.205 95.495 93.375 95.665 ;
        RECT 93.665 95.495 93.835 95.665 ;
        RECT 94.125 95.495 94.295 95.665 ;
        RECT 94.585 95.495 94.755 95.665 ;
        RECT 95.045 95.495 95.215 95.665 ;
        RECT 95.505 95.495 95.675 95.665 ;
        RECT 95.965 95.495 96.135 95.665 ;
        RECT 96.425 95.495 96.595 95.665 ;
        RECT 96.885 95.495 97.055 95.665 ;
        RECT 97.345 95.495 97.515 95.665 ;
        RECT 97.805 95.495 97.975 95.665 ;
        RECT 98.265 95.495 98.435 95.665 ;
        RECT 98.725 95.495 98.895 95.665 ;
        RECT 99.185 95.495 99.355 95.665 ;
        RECT 99.645 95.495 99.815 95.665 ;
        RECT 16.845 90.055 17.015 90.225 ;
        RECT 17.305 90.055 17.475 90.225 ;
        RECT 17.765 90.055 17.935 90.225 ;
        RECT 18.225 90.055 18.395 90.225 ;
        RECT 18.685 90.055 18.855 90.225 ;
        RECT 19.145 90.055 19.315 90.225 ;
        RECT 19.605 90.055 19.775 90.225 ;
        RECT 20.065 90.055 20.235 90.225 ;
        RECT 20.525 90.055 20.695 90.225 ;
        RECT 20.985 90.055 21.155 90.225 ;
        RECT 21.445 90.055 21.615 90.225 ;
        RECT 21.905 90.055 22.075 90.225 ;
        RECT 22.365 90.055 22.535 90.225 ;
        RECT 22.825 90.055 22.995 90.225 ;
        RECT 23.285 90.055 23.455 90.225 ;
        RECT 23.745 90.055 23.915 90.225 ;
        RECT 24.205 90.055 24.375 90.225 ;
        RECT 24.665 90.055 24.835 90.225 ;
        RECT 25.125 90.055 25.295 90.225 ;
        RECT 25.585 90.055 25.755 90.225 ;
        RECT 26.045 90.055 26.215 90.225 ;
        RECT 26.505 90.055 26.675 90.225 ;
        RECT 26.965 90.055 27.135 90.225 ;
        RECT 27.425 90.055 27.595 90.225 ;
        RECT 27.885 90.055 28.055 90.225 ;
        RECT 28.345 90.055 28.515 90.225 ;
        RECT 28.805 90.055 28.975 90.225 ;
        RECT 29.265 90.055 29.435 90.225 ;
        RECT 29.725 90.055 29.895 90.225 ;
        RECT 30.185 90.055 30.355 90.225 ;
        RECT 30.645 90.055 30.815 90.225 ;
        RECT 31.105 90.055 31.275 90.225 ;
        RECT 31.565 90.055 31.735 90.225 ;
        RECT 32.025 90.055 32.195 90.225 ;
        RECT 32.485 90.055 32.655 90.225 ;
        RECT 32.945 90.055 33.115 90.225 ;
        RECT 33.405 90.055 33.575 90.225 ;
        RECT 33.865 90.055 34.035 90.225 ;
        RECT 34.325 90.055 34.495 90.225 ;
        RECT 34.785 90.055 34.955 90.225 ;
        RECT 35.245 90.055 35.415 90.225 ;
        RECT 35.705 90.055 35.875 90.225 ;
        RECT 36.165 90.055 36.335 90.225 ;
        RECT 36.625 90.055 36.795 90.225 ;
        RECT 37.085 90.055 37.255 90.225 ;
        RECT 37.545 90.055 37.715 90.225 ;
        RECT 38.005 90.055 38.175 90.225 ;
        RECT 38.465 90.055 38.635 90.225 ;
        RECT 38.925 90.055 39.095 90.225 ;
        RECT 39.385 90.055 39.555 90.225 ;
        RECT 39.845 90.055 40.015 90.225 ;
        RECT 40.305 90.055 40.475 90.225 ;
        RECT 40.765 90.055 40.935 90.225 ;
        RECT 41.225 90.055 41.395 90.225 ;
        RECT 41.685 90.055 41.855 90.225 ;
        RECT 42.145 90.055 42.315 90.225 ;
        RECT 42.605 90.055 42.775 90.225 ;
        RECT 43.065 90.055 43.235 90.225 ;
        RECT 43.525 90.055 43.695 90.225 ;
        RECT 43.985 90.055 44.155 90.225 ;
        RECT 44.445 90.055 44.615 90.225 ;
        RECT 44.905 90.055 45.075 90.225 ;
        RECT 45.365 90.055 45.535 90.225 ;
        RECT 45.825 90.055 45.995 90.225 ;
        RECT 46.285 90.055 46.455 90.225 ;
        RECT 46.745 90.055 46.915 90.225 ;
        RECT 47.205 90.055 47.375 90.225 ;
        RECT 47.665 90.055 47.835 90.225 ;
        RECT 48.125 90.055 48.295 90.225 ;
        RECT 48.585 90.055 48.755 90.225 ;
        RECT 49.045 90.055 49.215 90.225 ;
        RECT 49.505 90.055 49.675 90.225 ;
        RECT 49.965 90.055 50.135 90.225 ;
        RECT 50.425 90.055 50.595 90.225 ;
        RECT 50.885 90.055 51.055 90.225 ;
        RECT 51.345 90.055 51.515 90.225 ;
        RECT 51.805 90.055 51.975 90.225 ;
        RECT 52.265 90.055 52.435 90.225 ;
        RECT 52.725 90.055 52.895 90.225 ;
        RECT 53.185 90.055 53.355 90.225 ;
        RECT 53.645 90.055 53.815 90.225 ;
        RECT 54.105 90.055 54.275 90.225 ;
        RECT 54.565 90.055 54.735 90.225 ;
        RECT 55.025 90.055 55.195 90.225 ;
        RECT 55.485 90.055 55.655 90.225 ;
        RECT 55.945 90.055 56.115 90.225 ;
        RECT 56.405 90.055 56.575 90.225 ;
        RECT 56.865 90.055 57.035 90.225 ;
        RECT 57.325 90.055 57.495 90.225 ;
        RECT 57.785 90.055 57.955 90.225 ;
        RECT 58.245 90.055 58.415 90.225 ;
        RECT 58.705 90.055 58.875 90.225 ;
        RECT 59.165 90.055 59.335 90.225 ;
        RECT 59.625 90.055 59.795 90.225 ;
        RECT 60.085 90.055 60.255 90.225 ;
        RECT 60.545 90.055 60.715 90.225 ;
        RECT 61.005 90.055 61.175 90.225 ;
        RECT 61.465 90.055 61.635 90.225 ;
        RECT 61.925 90.055 62.095 90.225 ;
        RECT 62.385 90.055 62.555 90.225 ;
        RECT 62.845 90.055 63.015 90.225 ;
        RECT 63.305 90.055 63.475 90.225 ;
        RECT 63.765 90.055 63.935 90.225 ;
        RECT 64.225 90.055 64.395 90.225 ;
        RECT 64.685 90.055 64.855 90.225 ;
        RECT 65.145 90.055 65.315 90.225 ;
        RECT 65.605 90.055 65.775 90.225 ;
        RECT 66.065 90.055 66.235 90.225 ;
        RECT 66.525 90.055 66.695 90.225 ;
        RECT 66.985 90.055 67.155 90.225 ;
        RECT 67.445 90.055 67.615 90.225 ;
        RECT 67.905 90.055 68.075 90.225 ;
        RECT 68.365 90.055 68.535 90.225 ;
        RECT 68.825 90.055 68.995 90.225 ;
        RECT 69.285 90.055 69.455 90.225 ;
        RECT 69.745 90.055 69.915 90.225 ;
        RECT 70.205 90.055 70.375 90.225 ;
        RECT 70.665 90.055 70.835 90.225 ;
        RECT 71.125 90.055 71.295 90.225 ;
        RECT 71.585 90.055 71.755 90.225 ;
        RECT 72.045 90.055 72.215 90.225 ;
        RECT 72.505 90.055 72.675 90.225 ;
        RECT 72.965 90.055 73.135 90.225 ;
        RECT 73.425 90.055 73.595 90.225 ;
        RECT 73.885 90.055 74.055 90.225 ;
        RECT 74.345 90.055 74.515 90.225 ;
        RECT 74.805 90.055 74.975 90.225 ;
        RECT 75.265 90.055 75.435 90.225 ;
        RECT 75.725 90.055 75.895 90.225 ;
        RECT 76.185 90.055 76.355 90.225 ;
        RECT 76.645 90.055 76.815 90.225 ;
        RECT 77.105 90.055 77.275 90.225 ;
        RECT 77.565 90.055 77.735 90.225 ;
        RECT 78.025 90.055 78.195 90.225 ;
        RECT 78.485 90.055 78.655 90.225 ;
        RECT 78.945 90.055 79.115 90.225 ;
        RECT 79.405 90.055 79.575 90.225 ;
        RECT 79.865 90.055 80.035 90.225 ;
        RECT 80.325 90.055 80.495 90.225 ;
        RECT 80.785 90.055 80.955 90.225 ;
        RECT 81.245 90.055 81.415 90.225 ;
        RECT 81.705 90.055 81.875 90.225 ;
        RECT 82.165 90.055 82.335 90.225 ;
        RECT 82.625 90.055 82.795 90.225 ;
        RECT 83.085 90.055 83.255 90.225 ;
        RECT 83.545 90.055 83.715 90.225 ;
        RECT 84.005 90.055 84.175 90.225 ;
        RECT 84.465 90.055 84.635 90.225 ;
        RECT 84.925 90.055 85.095 90.225 ;
        RECT 85.385 90.055 85.555 90.225 ;
        RECT 85.845 90.055 86.015 90.225 ;
        RECT 86.305 90.055 86.475 90.225 ;
        RECT 86.765 90.055 86.935 90.225 ;
        RECT 87.225 90.055 87.395 90.225 ;
        RECT 87.685 90.055 87.855 90.225 ;
        RECT 88.145 90.055 88.315 90.225 ;
        RECT 88.605 90.055 88.775 90.225 ;
        RECT 89.065 90.055 89.235 90.225 ;
        RECT 89.525 90.055 89.695 90.225 ;
        RECT 89.985 90.055 90.155 90.225 ;
        RECT 90.445 90.055 90.615 90.225 ;
        RECT 90.905 90.055 91.075 90.225 ;
        RECT 91.365 90.055 91.535 90.225 ;
        RECT 91.825 90.055 91.995 90.225 ;
        RECT 92.285 90.055 92.455 90.225 ;
        RECT 92.745 90.055 92.915 90.225 ;
        RECT 93.205 90.055 93.375 90.225 ;
        RECT 93.665 90.055 93.835 90.225 ;
        RECT 94.125 90.055 94.295 90.225 ;
        RECT 94.585 90.055 94.755 90.225 ;
        RECT 95.045 90.055 95.215 90.225 ;
        RECT 95.505 90.055 95.675 90.225 ;
        RECT 95.965 90.055 96.135 90.225 ;
        RECT 96.425 90.055 96.595 90.225 ;
        RECT 96.885 90.055 97.055 90.225 ;
        RECT 97.345 90.055 97.515 90.225 ;
        RECT 97.805 90.055 97.975 90.225 ;
        RECT 98.265 90.055 98.435 90.225 ;
        RECT 98.725 90.055 98.895 90.225 ;
        RECT 99.185 90.055 99.355 90.225 ;
        RECT 99.645 90.055 99.815 90.225 ;
        RECT 16.845 84.615 17.015 84.785 ;
        RECT 17.305 84.615 17.475 84.785 ;
        RECT 17.765 84.615 17.935 84.785 ;
        RECT 18.225 84.615 18.395 84.785 ;
        RECT 18.685 84.615 18.855 84.785 ;
        RECT 19.145 84.615 19.315 84.785 ;
        RECT 19.605 84.615 19.775 84.785 ;
        RECT 20.065 84.615 20.235 84.785 ;
        RECT 20.525 84.615 20.695 84.785 ;
        RECT 20.985 84.615 21.155 84.785 ;
        RECT 21.445 84.615 21.615 84.785 ;
        RECT 21.905 84.615 22.075 84.785 ;
        RECT 22.365 84.615 22.535 84.785 ;
        RECT 22.825 84.615 22.995 84.785 ;
        RECT 23.285 84.615 23.455 84.785 ;
        RECT 23.745 84.615 23.915 84.785 ;
        RECT 24.205 84.615 24.375 84.785 ;
        RECT 24.665 84.615 24.835 84.785 ;
        RECT 25.125 84.615 25.295 84.785 ;
        RECT 25.585 84.615 25.755 84.785 ;
        RECT 26.045 84.615 26.215 84.785 ;
        RECT 26.505 84.615 26.675 84.785 ;
        RECT 26.965 84.615 27.135 84.785 ;
        RECT 27.425 84.615 27.595 84.785 ;
        RECT 27.885 84.615 28.055 84.785 ;
        RECT 28.345 84.615 28.515 84.785 ;
        RECT 28.805 84.615 28.975 84.785 ;
        RECT 29.265 84.615 29.435 84.785 ;
        RECT 29.725 84.615 29.895 84.785 ;
        RECT 30.185 84.615 30.355 84.785 ;
        RECT 30.645 84.615 30.815 84.785 ;
        RECT 31.105 84.615 31.275 84.785 ;
        RECT 31.565 84.615 31.735 84.785 ;
        RECT 32.025 84.615 32.195 84.785 ;
        RECT 32.485 84.615 32.655 84.785 ;
        RECT 32.945 84.615 33.115 84.785 ;
        RECT 33.405 84.615 33.575 84.785 ;
        RECT 33.865 84.615 34.035 84.785 ;
        RECT 34.325 84.615 34.495 84.785 ;
        RECT 34.785 84.615 34.955 84.785 ;
        RECT 35.245 84.615 35.415 84.785 ;
        RECT 35.705 84.615 35.875 84.785 ;
        RECT 36.165 84.615 36.335 84.785 ;
        RECT 36.625 84.615 36.795 84.785 ;
        RECT 37.085 84.615 37.255 84.785 ;
        RECT 37.545 84.615 37.715 84.785 ;
        RECT 38.005 84.615 38.175 84.785 ;
        RECT 38.465 84.615 38.635 84.785 ;
        RECT 38.925 84.615 39.095 84.785 ;
        RECT 39.385 84.615 39.555 84.785 ;
        RECT 39.845 84.615 40.015 84.785 ;
        RECT 40.305 84.615 40.475 84.785 ;
        RECT 40.765 84.615 40.935 84.785 ;
        RECT 41.225 84.615 41.395 84.785 ;
        RECT 41.685 84.615 41.855 84.785 ;
        RECT 42.145 84.615 42.315 84.785 ;
        RECT 42.605 84.615 42.775 84.785 ;
        RECT 43.065 84.615 43.235 84.785 ;
        RECT 43.525 84.615 43.695 84.785 ;
        RECT 43.985 84.615 44.155 84.785 ;
        RECT 44.445 84.615 44.615 84.785 ;
        RECT 44.905 84.615 45.075 84.785 ;
        RECT 45.365 84.615 45.535 84.785 ;
        RECT 45.825 84.615 45.995 84.785 ;
        RECT 46.285 84.615 46.455 84.785 ;
        RECT 46.745 84.615 46.915 84.785 ;
        RECT 47.205 84.615 47.375 84.785 ;
        RECT 47.665 84.615 47.835 84.785 ;
        RECT 48.125 84.615 48.295 84.785 ;
        RECT 48.585 84.615 48.755 84.785 ;
        RECT 49.045 84.615 49.215 84.785 ;
        RECT 49.505 84.615 49.675 84.785 ;
        RECT 49.965 84.615 50.135 84.785 ;
        RECT 50.425 84.615 50.595 84.785 ;
        RECT 50.885 84.615 51.055 84.785 ;
        RECT 51.345 84.615 51.515 84.785 ;
        RECT 51.805 84.615 51.975 84.785 ;
        RECT 52.265 84.615 52.435 84.785 ;
        RECT 52.725 84.615 52.895 84.785 ;
        RECT 53.185 84.615 53.355 84.785 ;
        RECT 53.645 84.615 53.815 84.785 ;
        RECT 54.105 84.615 54.275 84.785 ;
        RECT 54.565 84.615 54.735 84.785 ;
        RECT 55.025 84.615 55.195 84.785 ;
        RECT 55.485 84.615 55.655 84.785 ;
        RECT 55.945 84.615 56.115 84.785 ;
        RECT 56.405 84.615 56.575 84.785 ;
        RECT 56.865 84.615 57.035 84.785 ;
        RECT 57.325 84.615 57.495 84.785 ;
        RECT 57.785 84.615 57.955 84.785 ;
        RECT 58.245 84.615 58.415 84.785 ;
        RECT 58.705 84.615 58.875 84.785 ;
        RECT 59.165 84.615 59.335 84.785 ;
        RECT 59.625 84.615 59.795 84.785 ;
        RECT 60.085 84.615 60.255 84.785 ;
        RECT 60.545 84.615 60.715 84.785 ;
        RECT 61.005 84.615 61.175 84.785 ;
        RECT 61.465 84.615 61.635 84.785 ;
        RECT 61.925 84.615 62.095 84.785 ;
        RECT 62.385 84.615 62.555 84.785 ;
        RECT 62.845 84.615 63.015 84.785 ;
        RECT 63.305 84.615 63.475 84.785 ;
        RECT 63.765 84.615 63.935 84.785 ;
        RECT 64.225 84.615 64.395 84.785 ;
        RECT 64.685 84.615 64.855 84.785 ;
        RECT 65.145 84.615 65.315 84.785 ;
        RECT 65.605 84.615 65.775 84.785 ;
        RECT 66.065 84.615 66.235 84.785 ;
        RECT 66.525 84.615 66.695 84.785 ;
        RECT 66.985 84.615 67.155 84.785 ;
        RECT 67.445 84.615 67.615 84.785 ;
        RECT 67.905 84.615 68.075 84.785 ;
        RECT 68.365 84.615 68.535 84.785 ;
        RECT 68.825 84.615 68.995 84.785 ;
        RECT 69.285 84.615 69.455 84.785 ;
        RECT 69.745 84.615 69.915 84.785 ;
        RECT 70.205 84.615 70.375 84.785 ;
        RECT 70.665 84.615 70.835 84.785 ;
        RECT 71.125 84.615 71.295 84.785 ;
        RECT 71.585 84.615 71.755 84.785 ;
        RECT 72.045 84.615 72.215 84.785 ;
        RECT 72.505 84.615 72.675 84.785 ;
        RECT 72.965 84.615 73.135 84.785 ;
        RECT 73.425 84.615 73.595 84.785 ;
        RECT 73.885 84.615 74.055 84.785 ;
        RECT 74.345 84.615 74.515 84.785 ;
        RECT 74.805 84.615 74.975 84.785 ;
        RECT 75.265 84.615 75.435 84.785 ;
        RECT 75.725 84.615 75.895 84.785 ;
        RECT 76.185 84.615 76.355 84.785 ;
        RECT 76.645 84.615 76.815 84.785 ;
        RECT 77.105 84.615 77.275 84.785 ;
        RECT 77.565 84.615 77.735 84.785 ;
        RECT 78.025 84.615 78.195 84.785 ;
        RECT 78.485 84.615 78.655 84.785 ;
        RECT 78.945 84.615 79.115 84.785 ;
        RECT 79.405 84.615 79.575 84.785 ;
        RECT 79.865 84.615 80.035 84.785 ;
        RECT 80.325 84.615 80.495 84.785 ;
        RECT 80.785 84.615 80.955 84.785 ;
        RECT 81.245 84.615 81.415 84.785 ;
        RECT 81.705 84.615 81.875 84.785 ;
        RECT 82.165 84.615 82.335 84.785 ;
        RECT 82.625 84.615 82.795 84.785 ;
        RECT 83.085 84.615 83.255 84.785 ;
        RECT 83.545 84.615 83.715 84.785 ;
        RECT 84.005 84.615 84.175 84.785 ;
        RECT 84.465 84.615 84.635 84.785 ;
        RECT 84.925 84.615 85.095 84.785 ;
        RECT 85.385 84.615 85.555 84.785 ;
        RECT 85.845 84.615 86.015 84.785 ;
        RECT 86.305 84.615 86.475 84.785 ;
        RECT 86.765 84.615 86.935 84.785 ;
        RECT 87.225 84.615 87.395 84.785 ;
        RECT 87.685 84.615 87.855 84.785 ;
        RECT 88.145 84.615 88.315 84.785 ;
        RECT 88.605 84.615 88.775 84.785 ;
        RECT 89.065 84.615 89.235 84.785 ;
        RECT 89.525 84.615 89.695 84.785 ;
        RECT 89.985 84.615 90.155 84.785 ;
        RECT 90.445 84.615 90.615 84.785 ;
        RECT 90.905 84.615 91.075 84.785 ;
        RECT 91.365 84.615 91.535 84.785 ;
        RECT 91.825 84.615 91.995 84.785 ;
        RECT 92.285 84.615 92.455 84.785 ;
        RECT 92.745 84.615 92.915 84.785 ;
        RECT 93.205 84.615 93.375 84.785 ;
        RECT 93.665 84.615 93.835 84.785 ;
        RECT 94.125 84.615 94.295 84.785 ;
        RECT 94.585 84.615 94.755 84.785 ;
        RECT 95.045 84.615 95.215 84.785 ;
        RECT 95.505 84.615 95.675 84.785 ;
        RECT 95.965 84.615 96.135 84.785 ;
        RECT 96.425 84.615 96.595 84.785 ;
        RECT 96.885 84.615 97.055 84.785 ;
        RECT 97.345 84.615 97.515 84.785 ;
        RECT 97.805 84.615 97.975 84.785 ;
        RECT 98.265 84.615 98.435 84.785 ;
        RECT 98.725 84.615 98.895 84.785 ;
        RECT 99.185 84.615 99.355 84.785 ;
        RECT 99.645 84.615 99.815 84.785 ;
        RECT 16.845 79.175 17.015 79.345 ;
        RECT 17.305 79.175 17.475 79.345 ;
        RECT 17.765 79.175 17.935 79.345 ;
        RECT 18.225 79.175 18.395 79.345 ;
        RECT 18.685 79.175 18.855 79.345 ;
        RECT 19.145 79.175 19.315 79.345 ;
        RECT 19.605 79.175 19.775 79.345 ;
        RECT 20.065 79.175 20.235 79.345 ;
        RECT 20.525 79.175 20.695 79.345 ;
        RECT 20.985 79.175 21.155 79.345 ;
        RECT 21.445 79.175 21.615 79.345 ;
        RECT 21.905 79.175 22.075 79.345 ;
        RECT 22.365 79.175 22.535 79.345 ;
        RECT 22.825 79.175 22.995 79.345 ;
        RECT 23.285 79.175 23.455 79.345 ;
        RECT 23.745 79.175 23.915 79.345 ;
        RECT 24.205 79.175 24.375 79.345 ;
        RECT 24.665 79.175 24.835 79.345 ;
        RECT 25.125 79.175 25.295 79.345 ;
        RECT 25.585 79.175 25.755 79.345 ;
        RECT 26.045 79.175 26.215 79.345 ;
        RECT 26.505 79.175 26.675 79.345 ;
        RECT 26.965 79.175 27.135 79.345 ;
        RECT 27.425 79.175 27.595 79.345 ;
        RECT 27.885 79.175 28.055 79.345 ;
        RECT 28.345 79.175 28.515 79.345 ;
        RECT 28.805 79.175 28.975 79.345 ;
        RECT 29.265 79.175 29.435 79.345 ;
        RECT 29.725 79.175 29.895 79.345 ;
        RECT 30.185 79.175 30.355 79.345 ;
        RECT 30.645 79.175 30.815 79.345 ;
        RECT 31.105 79.175 31.275 79.345 ;
        RECT 31.565 79.175 31.735 79.345 ;
        RECT 32.025 79.175 32.195 79.345 ;
        RECT 32.485 79.175 32.655 79.345 ;
        RECT 32.945 79.175 33.115 79.345 ;
        RECT 33.405 79.175 33.575 79.345 ;
        RECT 33.865 79.175 34.035 79.345 ;
        RECT 34.325 79.175 34.495 79.345 ;
        RECT 34.785 79.175 34.955 79.345 ;
        RECT 35.245 79.175 35.415 79.345 ;
        RECT 35.705 79.175 35.875 79.345 ;
        RECT 36.165 79.175 36.335 79.345 ;
        RECT 36.625 79.175 36.795 79.345 ;
        RECT 37.085 79.175 37.255 79.345 ;
        RECT 37.545 79.175 37.715 79.345 ;
        RECT 38.005 79.175 38.175 79.345 ;
        RECT 38.465 79.175 38.635 79.345 ;
        RECT 38.925 79.175 39.095 79.345 ;
        RECT 39.385 79.175 39.555 79.345 ;
        RECT 39.845 79.175 40.015 79.345 ;
        RECT 40.305 79.175 40.475 79.345 ;
        RECT 40.765 79.175 40.935 79.345 ;
        RECT 41.225 79.175 41.395 79.345 ;
        RECT 41.685 79.175 41.855 79.345 ;
        RECT 42.145 79.175 42.315 79.345 ;
        RECT 42.605 79.175 42.775 79.345 ;
        RECT 43.065 79.175 43.235 79.345 ;
        RECT 43.525 79.175 43.695 79.345 ;
        RECT 43.985 79.175 44.155 79.345 ;
        RECT 44.445 79.175 44.615 79.345 ;
        RECT 44.905 79.175 45.075 79.345 ;
        RECT 45.365 79.175 45.535 79.345 ;
        RECT 45.825 79.175 45.995 79.345 ;
        RECT 46.285 79.175 46.455 79.345 ;
        RECT 46.745 79.175 46.915 79.345 ;
        RECT 47.205 79.175 47.375 79.345 ;
        RECT 47.665 79.175 47.835 79.345 ;
        RECT 48.125 79.175 48.295 79.345 ;
        RECT 48.585 79.175 48.755 79.345 ;
        RECT 49.045 79.175 49.215 79.345 ;
        RECT 49.505 79.175 49.675 79.345 ;
        RECT 49.965 79.175 50.135 79.345 ;
        RECT 50.425 79.175 50.595 79.345 ;
        RECT 50.885 79.175 51.055 79.345 ;
        RECT 51.345 79.175 51.515 79.345 ;
        RECT 51.805 79.175 51.975 79.345 ;
        RECT 52.265 79.175 52.435 79.345 ;
        RECT 52.725 79.175 52.895 79.345 ;
        RECT 53.185 79.175 53.355 79.345 ;
        RECT 53.645 79.175 53.815 79.345 ;
        RECT 54.105 79.175 54.275 79.345 ;
        RECT 54.565 79.175 54.735 79.345 ;
        RECT 55.025 79.175 55.195 79.345 ;
        RECT 55.485 79.175 55.655 79.345 ;
        RECT 55.945 79.175 56.115 79.345 ;
        RECT 56.405 79.175 56.575 79.345 ;
        RECT 56.865 79.175 57.035 79.345 ;
        RECT 57.325 79.175 57.495 79.345 ;
        RECT 57.785 79.175 57.955 79.345 ;
        RECT 58.245 79.175 58.415 79.345 ;
        RECT 58.705 79.175 58.875 79.345 ;
        RECT 59.165 79.175 59.335 79.345 ;
        RECT 59.625 79.175 59.795 79.345 ;
        RECT 60.085 79.175 60.255 79.345 ;
        RECT 60.545 79.175 60.715 79.345 ;
        RECT 61.005 79.175 61.175 79.345 ;
        RECT 61.465 79.175 61.635 79.345 ;
        RECT 61.925 79.175 62.095 79.345 ;
        RECT 62.385 79.175 62.555 79.345 ;
        RECT 62.845 79.175 63.015 79.345 ;
        RECT 63.305 79.175 63.475 79.345 ;
        RECT 63.765 79.175 63.935 79.345 ;
        RECT 64.225 79.175 64.395 79.345 ;
        RECT 64.685 79.175 64.855 79.345 ;
        RECT 65.145 79.175 65.315 79.345 ;
        RECT 65.605 79.175 65.775 79.345 ;
        RECT 66.065 79.175 66.235 79.345 ;
        RECT 66.525 79.175 66.695 79.345 ;
        RECT 66.985 79.175 67.155 79.345 ;
        RECT 67.445 79.175 67.615 79.345 ;
        RECT 67.905 79.175 68.075 79.345 ;
        RECT 68.365 79.175 68.535 79.345 ;
        RECT 68.825 79.175 68.995 79.345 ;
        RECT 69.285 79.175 69.455 79.345 ;
        RECT 69.745 79.175 69.915 79.345 ;
        RECT 70.205 79.175 70.375 79.345 ;
        RECT 70.665 79.175 70.835 79.345 ;
        RECT 71.125 79.175 71.295 79.345 ;
        RECT 71.585 79.175 71.755 79.345 ;
        RECT 72.045 79.175 72.215 79.345 ;
        RECT 72.505 79.175 72.675 79.345 ;
        RECT 72.965 79.175 73.135 79.345 ;
        RECT 73.425 79.175 73.595 79.345 ;
        RECT 73.885 79.175 74.055 79.345 ;
        RECT 74.345 79.175 74.515 79.345 ;
        RECT 74.805 79.175 74.975 79.345 ;
        RECT 75.265 79.175 75.435 79.345 ;
        RECT 75.725 79.175 75.895 79.345 ;
        RECT 76.185 79.175 76.355 79.345 ;
        RECT 76.645 79.175 76.815 79.345 ;
        RECT 77.105 79.175 77.275 79.345 ;
        RECT 77.565 79.175 77.735 79.345 ;
        RECT 78.025 79.175 78.195 79.345 ;
        RECT 78.485 79.175 78.655 79.345 ;
        RECT 78.945 79.175 79.115 79.345 ;
        RECT 79.405 79.175 79.575 79.345 ;
        RECT 79.865 79.175 80.035 79.345 ;
        RECT 80.325 79.175 80.495 79.345 ;
        RECT 80.785 79.175 80.955 79.345 ;
        RECT 81.245 79.175 81.415 79.345 ;
        RECT 81.705 79.175 81.875 79.345 ;
        RECT 82.165 79.175 82.335 79.345 ;
        RECT 82.625 79.175 82.795 79.345 ;
        RECT 83.085 79.175 83.255 79.345 ;
        RECT 83.545 79.175 83.715 79.345 ;
        RECT 84.005 79.175 84.175 79.345 ;
        RECT 84.465 79.175 84.635 79.345 ;
        RECT 84.925 79.175 85.095 79.345 ;
        RECT 85.385 79.175 85.555 79.345 ;
        RECT 85.845 79.175 86.015 79.345 ;
        RECT 86.305 79.175 86.475 79.345 ;
        RECT 86.765 79.175 86.935 79.345 ;
        RECT 87.225 79.175 87.395 79.345 ;
        RECT 87.685 79.175 87.855 79.345 ;
        RECT 88.145 79.175 88.315 79.345 ;
        RECT 88.605 79.175 88.775 79.345 ;
        RECT 89.065 79.175 89.235 79.345 ;
        RECT 89.525 79.175 89.695 79.345 ;
        RECT 89.985 79.175 90.155 79.345 ;
        RECT 90.445 79.175 90.615 79.345 ;
        RECT 90.905 79.175 91.075 79.345 ;
        RECT 91.365 79.175 91.535 79.345 ;
        RECT 91.825 79.175 91.995 79.345 ;
        RECT 92.285 79.175 92.455 79.345 ;
        RECT 92.745 79.175 92.915 79.345 ;
        RECT 93.205 79.175 93.375 79.345 ;
        RECT 93.665 79.175 93.835 79.345 ;
        RECT 94.125 79.175 94.295 79.345 ;
        RECT 94.585 79.175 94.755 79.345 ;
        RECT 95.045 79.175 95.215 79.345 ;
        RECT 95.505 79.175 95.675 79.345 ;
        RECT 95.965 79.175 96.135 79.345 ;
        RECT 96.425 79.175 96.595 79.345 ;
        RECT 96.885 79.175 97.055 79.345 ;
        RECT 97.345 79.175 97.515 79.345 ;
        RECT 97.805 79.175 97.975 79.345 ;
        RECT 98.265 79.175 98.435 79.345 ;
        RECT 98.725 79.175 98.895 79.345 ;
        RECT 99.185 79.175 99.355 79.345 ;
        RECT 99.645 79.175 99.815 79.345 ;
        RECT 16.845 73.735 17.015 73.905 ;
        RECT 17.305 73.735 17.475 73.905 ;
        RECT 17.765 73.735 17.935 73.905 ;
        RECT 18.225 73.735 18.395 73.905 ;
        RECT 18.685 73.735 18.855 73.905 ;
        RECT 19.145 73.735 19.315 73.905 ;
        RECT 19.605 73.735 19.775 73.905 ;
        RECT 20.065 73.735 20.235 73.905 ;
        RECT 20.525 73.735 20.695 73.905 ;
        RECT 20.985 73.735 21.155 73.905 ;
        RECT 21.445 73.735 21.615 73.905 ;
        RECT 21.905 73.735 22.075 73.905 ;
        RECT 22.365 73.735 22.535 73.905 ;
        RECT 22.825 73.735 22.995 73.905 ;
        RECT 23.285 73.735 23.455 73.905 ;
        RECT 23.745 73.735 23.915 73.905 ;
        RECT 24.205 73.735 24.375 73.905 ;
        RECT 24.665 73.735 24.835 73.905 ;
        RECT 25.125 73.735 25.295 73.905 ;
        RECT 25.585 73.735 25.755 73.905 ;
        RECT 26.045 73.735 26.215 73.905 ;
        RECT 26.505 73.735 26.675 73.905 ;
        RECT 26.965 73.735 27.135 73.905 ;
        RECT 27.425 73.735 27.595 73.905 ;
        RECT 27.885 73.735 28.055 73.905 ;
        RECT 28.345 73.735 28.515 73.905 ;
        RECT 28.805 73.735 28.975 73.905 ;
        RECT 29.265 73.735 29.435 73.905 ;
        RECT 29.725 73.735 29.895 73.905 ;
        RECT 30.185 73.735 30.355 73.905 ;
        RECT 30.645 73.735 30.815 73.905 ;
        RECT 31.105 73.735 31.275 73.905 ;
        RECT 31.565 73.735 31.735 73.905 ;
        RECT 32.025 73.735 32.195 73.905 ;
        RECT 32.485 73.735 32.655 73.905 ;
        RECT 32.945 73.735 33.115 73.905 ;
        RECT 33.405 73.735 33.575 73.905 ;
        RECT 33.865 73.735 34.035 73.905 ;
        RECT 34.325 73.735 34.495 73.905 ;
        RECT 34.785 73.735 34.955 73.905 ;
        RECT 35.245 73.735 35.415 73.905 ;
        RECT 35.705 73.735 35.875 73.905 ;
        RECT 36.165 73.735 36.335 73.905 ;
        RECT 36.625 73.735 36.795 73.905 ;
        RECT 37.085 73.735 37.255 73.905 ;
        RECT 37.545 73.735 37.715 73.905 ;
        RECT 38.005 73.735 38.175 73.905 ;
        RECT 38.465 73.735 38.635 73.905 ;
        RECT 38.925 73.735 39.095 73.905 ;
        RECT 39.385 73.735 39.555 73.905 ;
        RECT 39.845 73.735 40.015 73.905 ;
        RECT 40.305 73.735 40.475 73.905 ;
        RECT 40.765 73.735 40.935 73.905 ;
        RECT 41.225 73.735 41.395 73.905 ;
        RECT 41.685 73.735 41.855 73.905 ;
        RECT 42.145 73.735 42.315 73.905 ;
        RECT 42.605 73.735 42.775 73.905 ;
        RECT 43.065 73.735 43.235 73.905 ;
        RECT 43.525 73.735 43.695 73.905 ;
        RECT 43.985 73.735 44.155 73.905 ;
        RECT 44.445 73.735 44.615 73.905 ;
        RECT 44.905 73.735 45.075 73.905 ;
        RECT 45.365 73.735 45.535 73.905 ;
        RECT 45.825 73.735 45.995 73.905 ;
        RECT 46.285 73.735 46.455 73.905 ;
        RECT 46.745 73.735 46.915 73.905 ;
        RECT 47.205 73.735 47.375 73.905 ;
        RECT 47.665 73.735 47.835 73.905 ;
        RECT 48.125 73.735 48.295 73.905 ;
        RECT 48.585 73.735 48.755 73.905 ;
        RECT 49.045 73.735 49.215 73.905 ;
        RECT 49.505 73.735 49.675 73.905 ;
        RECT 49.965 73.735 50.135 73.905 ;
        RECT 50.425 73.735 50.595 73.905 ;
        RECT 50.885 73.735 51.055 73.905 ;
        RECT 51.345 73.735 51.515 73.905 ;
        RECT 51.805 73.735 51.975 73.905 ;
        RECT 52.265 73.735 52.435 73.905 ;
        RECT 52.725 73.735 52.895 73.905 ;
        RECT 53.185 73.735 53.355 73.905 ;
        RECT 53.645 73.735 53.815 73.905 ;
        RECT 54.105 73.735 54.275 73.905 ;
        RECT 54.565 73.735 54.735 73.905 ;
        RECT 55.025 73.735 55.195 73.905 ;
        RECT 55.485 73.735 55.655 73.905 ;
        RECT 55.945 73.735 56.115 73.905 ;
        RECT 56.405 73.735 56.575 73.905 ;
        RECT 56.865 73.735 57.035 73.905 ;
        RECT 57.325 73.735 57.495 73.905 ;
        RECT 57.785 73.735 57.955 73.905 ;
        RECT 58.245 73.735 58.415 73.905 ;
        RECT 58.705 73.735 58.875 73.905 ;
        RECT 59.165 73.735 59.335 73.905 ;
        RECT 59.625 73.735 59.795 73.905 ;
        RECT 60.085 73.735 60.255 73.905 ;
        RECT 60.545 73.735 60.715 73.905 ;
        RECT 61.005 73.735 61.175 73.905 ;
        RECT 61.465 73.735 61.635 73.905 ;
        RECT 61.925 73.735 62.095 73.905 ;
        RECT 62.385 73.735 62.555 73.905 ;
        RECT 62.845 73.735 63.015 73.905 ;
        RECT 63.305 73.735 63.475 73.905 ;
        RECT 63.765 73.735 63.935 73.905 ;
        RECT 64.225 73.735 64.395 73.905 ;
        RECT 64.685 73.735 64.855 73.905 ;
        RECT 65.145 73.735 65.315 73.905 ;
        RECT 65.605 73.735 65.775 73.905 ;
        RECT 66.065 73.735 66.235 73.905 ;
        RECT 66.525 73.735 66.695 73.905 ;
        RECT 66.985 73.735 67.155 73.905 ;
        RECT 67.445 73.735 67.615 73.905 ;
        RECT 67.905 73.735 68.075 73.905 ;
        RECT 68.365 73.735 68.535 73.905 ;
        RECT 68.825 73.735 68.995 73.905 ;
        RECT 69.285 73.735 69.455 73.905 ;
        RECT 69.745 73.735 69.915 73.905 ;
        RECT 70.205 73.735 70.375 73.905 ;
        RECT 70.665 73.735 70.835 73.905 ;
        RECT 71.125 73.735 71.295 73.905 ;
        RECT 71.585 73.735 71.755 73.905 ;
        RECT 72.045 73.735 72.215 73.905 ;
        RECT 72.505 73.735 72.675 73.905 ;
        RECT 72.965 73.735 73.135 73.905 ;
        RECT 73.425 73.735 73.595 73.905 ;
        RECT 73.885 73.735 74.055 73.905 ;
        RECT 74.345 73.735 74.515 73.905 ;
        RECT 74.805 73.735 74.975 73.905 ;
        RECT 75.265 73.735 75.435 73.905 ;
        RECT 75.725 73.735 75.895 73.905 ;
        RECT 76.185 73.735 76.355 73.905 ;
        RECT 76.645 73.735 76.815 73.905 ;
        RECT 77.105 73.735 77.275 73.905 ;
        RECT 77.565 73.735 77.735 73.905 ;
        RECT 78.025 73.735 78.195 73.905 ;
        RECT 78.485 73.735 78.655 73.905 ;
        RECT 78.945 73.735 79.115 73.905 ;
        RECT 79.405 73.735 79.575 73.905 ;
        RECT 79.865 73.735 80.035 73.905 ;
        RECT 80.325 73.735 80.495 73.905 ;
        RECT 80.785 73.735 80.955 73.905 ;
        RECT 81.245 73.735 81.415 73.905 ;
        RECT 81.705 73.735 81.875 73.905 ;
        RECT 82.165 73.735 82.335 73.905 ;
        RECT 82.625 73.735 82.795 73.905 ;
        RECT 83.085 73.735 83.255 73.905 ;
        RECT 83.545 73.735 83.715 73.905 ;
        RECT 84.005 73.735 84.175 73.905 ;
        RECT 84.465 73.735 84.635 73.905 ;
        RECT 84.925 73.735 85.095 73.905 ;
        RECT 85.385 73.735 85.555 73.905 ;
        RECT 85.845 73.735 86.015 73.905 ;
        RECT 86.305 73.735 86.475 73.905 ;
        RECT 86.765 73.735 86.935 73.905 ;
        RECT 87.225 73.735 87.395 73.905 ;
        RECT 87.685 73.735 87.855 73.905 ;
        RECT 88.145 73.735 88.315 73.905 ;
        RECT 88.605 73.735 88.775 73.905 ;
        RECT 89.065 73.735 89.235 73.905 ;
        RECT 89.525 73.735 89.695 73.905 ;
        RECT 89.985 73.735 90.155 73.905 ;
        RECT 90.445 73.735 90.615 73.905 ;
        RECT 90.905 73.735 91.075 73.905 ;
        RECT 91.365 73.735 91.535 73.905 ;
        RECT 91.825 73.735 91.995 73.905 ;
        RECT 92.285 73.735 92.455 73.905 ;
        RECT 92.745 73.735 92.915 73.905 ;
        RECT 93.205 73.735 93.375 73.905 ;
        RECT 93.665 73.735 93.835 73.905 ;
        RECT 94.125 73.735 94.295 73.905 ;
        RECT 94.585 73.735 94.755 73.905 ;
        RECT 95.045 73.735 95.215 73.905 ;
        RECT 95.505 73.735 95.675 73.905 ;
        RECT 95.965 73.735 96.135 73.905 ;
        RECT 96.425 73.735 96.595 73.905 ;
        RECT 96.885 73.735 97.055 73.905 ;
        RECT 97.345 73.735 97.515 73.905 ;
        RECT 97.805 73.735 97.975 73.905 ;
        RECT 98.265 73.735 98.435 73.905 ;
        RECT 98.725 73.735 98.895 73.905 ;
        RECT 99.185 73.735 99.355 73.905 ;
        RECT 99.645 73.735 99.815 73.905 ;
        RECT 16.845 68.295 17.015 68.465 ;
        RECT 17.305 68.295 17.475 68.465 ;
        RECT 17.765 68.295 17.935 68.465 ;
        RECT 18.225 68.295 18.395 68.465 ;
        RECT 18.685 68.295 18.855 68.465 ;
        RECT 19.145 68.295 19.315 68.465 ;
        RECT 19.605 68.295 19.775 68.465 ;
        RECT 20.065 68.295 20.235 68.465 ;
        RECT 20.525 68.295 20.695 68.465 ;
        RECT 20.985 68.295 21.155 68.465 ;
        RECT 21.445 68.295 21.615 68.465 ;
        RECT 21.905 68.295 22.075 68.465 ;
        RECT 22.365 68.295 22.535 68.465 ;
        RECT 22.825 68.295 22.995 68.465 ;
        RECT 23.285 68.295 23.455 68.465 ;
        RECT 23.745 68.295 23.915 68.465 ;
        RECT 24.205 68.295 24.375 68.465 ;
        RECT 24.665 68.295 24.835 68.465 ;
        RECT 25.125 68.295 25.295 68.465 ;
        RECT 25.585 68.295 25.755 68.465 ;
        RECT 26.045 68.295 26.215 68.465 ;
        RECT 26.505 68.295 26.675 68.465 ;
        RECT 26.965 68.295 27.135 68.465 ;
        RECT 27.425 68.295 27.595 68.465 ;
        RECT 27.885 68.295 28.055 68.465 ;
        RECT 28.345 68.295 28.515 68.465 ;
        RECT 28.805 68.295 28.975 68.465 ;
        RECT 29.265 68.295 29.435 68.465 ;
        RECT 29.725 68.295 29.895 68.465 ;
        RECT 30.185 68.295 30.355 68.465 ;
        RECT 30.645 68.295 30.815 68.465 ;
        RECT 31.105 68.295 31.275 68.465 ;
        RECT 31.565 68.295 31.735 68.465 ;
        RECT 32.025 68.295 32.195 68.465 ;
        RECT 32.485 68.295 32.655 68.465 ;
        RECT 32.945 68.295 33.115 68.465 ;
        RECT 33.405 68.295 33.575 68.465 ;
        RECT 33.865 68.295 34.035 68.465 ;
        RECT 34.325 68.295 34.495 68.465 ;
        RECT 34.785 68.295 34.955 68.465 ;
        RECT 35.245 68.295 35.415 68.465 ;
        RECT 35.705 68.295 35.875 68.465 ;
        RECT 36.165 68.295 36.335 68.465 ;
        RECT 36.625 68.295 36.795 68.465 ;
        RECT 37.085 68.295 37.255 68.465 ;
        RECT 37.545 68.295 37.715 68.465 ;
        RECT 38.005 68.295 38.175 68.465 ;
        RECT 38.465 68.295 38.635 68.465 ;
        RECT 38.925 68.295 39.095 68.465 ;
        RECT 39.385 68.295 39.555 68.465 ;
        RECT 39.845 68.295 40.015 68.465 ;
        RECT 40.305 68.295 40.475 68.465 ;
        RECT 40.765 68.295 40.935 68.465 ;
        RECT 41.225 68.295 41.395 68.465 ;
        RECT 41.685 68.295 41.855 68.465 ;
        RECT 42.145 68.295 42.315 68.465 ;
        RECT 42.605 68.295 42.775 68.465 ;
        RECT 43.065 68.295 43.235 68.465 ;
        RECT 43.525 68.295 43.695 68.465 ;
        RECT 43.985 68.295 44.155 68.465 ;
        RECT 44.445 68.295 44.615 68.465 ;
        RECT 44.905 68.295 45.075 68.465 ;
        RECT 45.365 68.295 45.535 68.465 ;
        RECT 45.825 68.295 45.995 68.465 ;
        RECT 46.285 68.295 46.455 68.465 ;
        RECT 46.745 68.295 46.915 68.465 ;
        RECT 47.205 68.295 47.375 68.465 ;
        RECT 47.665 68.295 47.835 68.465 ;
        RECT 48.125 68.295 48.295 68.465 ;
        RECT 48.585 68.295 48.755 68.465 ;
        RECT 49.045 68.295 49.215 68.465 ;
        RECT 49.505 68.295 49.675 68.465 ;
        RECT 49.965 68.295 50.135 68.465 ;
        RECT 50.425 68.295 50.595 68.465 ;
        RECT 50.885 68.295 51.055 68.465 ;
        RECT 51.345 68.295 51.515 68.465 ;
        RECT 51.805 68.295 51.975 68.465 ;
        RECT 52.265 68.295 52.435 68.465 ;
        RECT 52.725 68.295 52.895 68.465 ;
        RECT 53.185 68.295 53.355 68.465 ;
        RECT 53.645 68.295 53.815 68.465 ;
        RECT 54.105 68.295 54.275 68.465 ;
        RECT 54.565 68.295 54.735 68.465 ;
        RECT 55.025 68.295 55.195 68.465 ;
        RECT 55.485 68.295 55.655 68.465 ;
        RECT 55.945 68.295 56.115 68.465 ;
        RECT 56.405 68.295 56.575 68.465 ;
        RECT 56.865 68.295 57.035 68.465 ;
        RECT 57.325 68.295 57.495 68.465 ;
        RECT 57.785 68.295 57.955 68.465 ;
        RECT 58.245 68.295 58.415 68.465 ;
        RECT 58.705 68.295 58.875 68.465 ;
        RECT 59.165 68.295 59.335 68.465 ;
        RECT 59.625 68.295 59.795 68.465 ;
        RECT 60.085 68.295 60.255 68.465 ;
        RECT 60.545 68.295 60.715 68.465 ;
        RECT 61.005 68.295 61.175 68.465 ;
        RECT 61.465 68.295 61.635 68.465 ;
        RECT 61.925 68.295 62.095 68.465 ;
        RECT 62.385 68.295 62.555 68.465 ;
        RECT 62.845 68.295 63.015 68.465 ;
        RECT 63.305 68.295 63.475 68.465 ;
        RECT 63.765 68.295 63.935 68.465 ;
        RECT 64.225 68.295 64.395 68.465 ;
        RECT 64.685 68.295 64.855 68.465 ;
        RECT 65.145 68.295 65.315 68.465 ;
        RECT 65.605 68.295 65.775 68.465 ;
        RECT 66.065 68.295 66.235 68.465 ;
        RECT 66.525 68.295 66.695 68.465 ;
        RECT 66.985 68.295 67.155 68.465 ;
        RECT 67.445 68.295 67.615 68.465 ;
        RECT 67.905 68.295 68.075 68.465 ;
        RECT 68.365 68.295 68.535 68.465 ;
        RECT 68.825 68.295 68.995 68.465 ;
        RECT 69.285 68.295 69.455 68.465 ;
        RECT 69.745 68.295 69.915 68.465 ;
        RECT 70.205 68.295 70.375 68.465 ;
        RECT 70.665 68.295 70.835 68.465 ;
        RECT 71.125 68.295 71.295 68.465 ;
        RECT 71.585 68.295 71.755 68.465 ;
        RECT 72.045 68.295 72.215 68.465 ;
        RECT 72.505 68.295 72.675 68.465 ;
        RECT 72.965 68.295 73.135 68.465 ;
        RECT 73.425 68.295 73.595 68.465 ;
        RECT 73.885 68.295 74.055 68.465 ;
        RECT 74.345 68.295 74.515 68.465 ;
        RECT 74.805 68.295 74.975 68.465 ;
        RECT 75.265 68.295 75.435 68.465 ;
        RECT 75.725 68.295 75.895 68.465 ;
        RECT 76.185 68.295 76.355 68.465 ;
        RECT 76.645 68.295 76.815 68.465 ;
        RECT 77.105 68.295 77.275 68.465 ;
        RECT 77.565 68.295 77.735 68.465 ;
        RECT 78.025 68.295 78.195 68.465 ;
        RECT 78.485 68.295 78.655 68.465 ;
        RECT 78.945 68.295 79.115 68.465 ;
        RECT 79.405 68.295 79.575 68.465 ;
        RECT 79.865 68.295 80.035 68.465 ;
        RECT 80.325 68.295 80.495 68.465 ;
        RECT 80.785 68.295 80.955 68.465 ;
        RECT 81.245 68.295 81.415 68.465 ;
        RECT 81.705 68.295 81.875 68.465 ;
        RECT 82.165 68.295 82.335 68.465 ;
        RECT 82.625 68.295 82.795 68.465 ;
        RECT 83.085 68.295 83.255 68.465 ;
        RECT 83.545 68.295 83.715 68.465 ;
        RECT 84.005 68.295 84.175 68.465 ;
        RECT 84.465 68.295 84.635 68.465 ;
        RECT 84.925 68.295 85.095 68.465 ;
        RECT 85.385 68.295 85.555 68.465 ;
        RECT 85.845 68.295 86.015 68.465 ;
        RECT 86.305 68.295 86.475 68.465 ;
        RECT 86.765 68.295 86.935 68.465 ;
        RECT 87.225 68.295 87.395 68.465 ;
        RECT 87.685 68.295 87.855 68.465 ;
        RECT 88.145 68.295 88.315 68.465 ;
        RECT 88.605 68.295 88.775 68.465 ;
        RECT 89.065 68.295 89.235 68.465 ;
        RECT 89.525 68.295 89.695 68.465 ;
        RECT 89.985 68.295 90.155 68.465 ;
        RECT 90.445 68.295 90.615 68.465 ;
        RECT 90.905 68.295 91.075 68.465 ;
        RECT 91.365 68.295 91.535 68.465 ;
        RECT 91.825 68.295 91.995 68.465 ;
        RECT 92.285 68.295 92.455 68.465 ;
        RECT 92.745 68.295 92.915 68.465 ;
        RECT 93.205 68.295 93.375 68.465 ;
        RECT 93.665 68.295 93.835 68.465 ;
        RECT 94.125 68.295 94.295 68.465 ;
        RECT 94.585 68.295 94.755 68.465 ;
        RECT 95.045 68.295 95.215 68.465 ;
        RECT 95.505 68.295 95.675 68.465 ;
        RECT 95.965 68.295 96.135 68.465 ;
        RECT 96.425 68.295 96.595 68.465 ;
        RECT 96.885 68.295 97.055 68.465 ;
        RECT 97.345 68.295 97.515 68.465 ;
        RECT 97.805 68.295 97.975 68.465 ;
        RECT 98.265 68.295 98.435 68.465 ;
        RECT 98.725 68.295 98.895 68.465 ;
        RECT 99.185 68.295 99.355 68.465 ;
        RECT 99.645 68.295 99.815 68.465 ;
        RECT 16.845 62.855 17.015 63.025 ;
        RECT 17.305 62.855 17.475 63.025 ;
        RECT 17.765 62.855 17.935 63.025 ;
        RECT 18.225 62.855 18.395 63.025 ;
        RECT 18.685 62.855 18.855 63.025 ;
        RECT 19.145 62.855 19.315 63.025 ;
        RECT 19.605 62.855 19.775 63.025 ;
        RECT 20.065 62.855 20.235 63.025 ;
        RECT 20.525 62.855 20.695 63.025 ;
        RECT 20.985 62.855 21.155 63.025 ;
        RECT 21.445 62.855 21.615 63.025 ;
        RECT 21.905 62.855 22.075 63.025 ;
        RECT 22.365 62.855 22.535 63.025 ;
        RECT 22.825 62.855 22.995 63.025 ;
        RECT 23.285 62.855 23.455 63.025 ;
        RECT 23.745 62.855 23.915 63.025 ;
        RECT 24.205 62.855 24.375 63.025 ;
        RECT 24.665 62.855 24.835 63.025 ;
        RECT 25.125 62.855 25.295 63.025 ;
        RECT 25.585 62.855 25.755 63.025 ;
        RECT 26.045 62.855 26.215 63.025 ;
        RECT 26.505 62.855 26.675 63.025 ;
        RECT 26.965 62.855 27.135 63.025 ;
        RECT 27.425 62.855 27.595 63.025 ;
        RECT 27.885 62.855 28.055 63.025 ;
        RECT 28.345 62.855 28.515 63.025 ;
        RECT 28.805 62.855 28.975 63.025 ;
        RECT 29.265 62.855 29.435 63.025 ;
        RECT 29.725 62.855 29.895 63.025 ;
        RECT 30.185 62.855 30.355 63.025 ;
        RECT 30.645 62.855 30.815 63.025 ;
        RECT 31.105 62.855 31.275 63.025 ;
        RECT 31.565 62.855 31.735 63.025 ;
        RECT 32.025 62.855 32.195 63.025 ;
        RECT 32.485 62.855 32.655 63.025 ;
        RECT 32.945 62.855 33.115 63.025 ;
        RECT 33.405 62.855 33.575 63.025 ;
        RECT 33.865 62.855 34.035 63.025 ;
        RECT 34.325 62.855 34.495 63.025 ;
        RECT 34.785 62.855 34.955 63.025 ;
        RECT 35.245 62.855 35.415 63.025 ;
        RECT 35.705 62.855 35.875 63.025 ;
        RECT 36.165 62.855 36.335 63.025 ;
        RECT 36.625 62.855 36.795 63.025 ;
        RECT 37.085 62.855 37.255 63.025 ;
        RECT 37.545 62.855 37.715 63.025 ;
        RECT 38.005 62.855 38.175 63.025 ;
        RECT 38.465 62.855 38.635 63.025 ;
        RECT 38.925 62.855 39.095 63.025 ;
        RECT 39.385 62.855 39.555 63.025 ;
        RECT 39.845 62.855 40.015 63.025 ;
        RECT 40.305 62.855 40.475 63.025 ;
        RECT 40.765 62.855 40.935 63.025 ;
        RECT 41.225 62.855 41.395 63.025 ;
        RECT 41.685 62.855 41.855 63.025 ;
        RECT 42.145 62.855 42.315 63.025 ;
        RECT 42.605 62.855 42.775 63.025 ;
        RECT 43.065 62.855 43.235 63.025 ;
        RECT 43.525 62.855 43.695 63.025 ;
        RECT 43.985 62.855 44.155 63.025 ;
        RECT 44.445 62.855 44.615 63.025 ;
        RECT 44.905 62.855 45.075 63.025 ;
        RECT 45.365 62.855 45.535 63.025 ;
        RECT 45.825 62.855 45.995 63.025 ;
        RECT 46.285 62.855 46.455 63.025 ;
        RECT 46.745 62.855 46.915 63.025 ;
        RECT 47.205 62.855 47.375 63.025 ;
        RECT 47.665 62.855 47.835 63.025 ;
        RECT 48.125 62.855 48.295 63.025 ;
        RECT 48.585 62.855 48.755 63.025 ;
        RECT 49.045 62.855 49.215 63.025 ;
        RECT 49.505 62.855 49.675 63.025 ;
        RECT 49.965 62.855 50.135 63.025 ;
        RECT 50.425 62.855 50.595 63.025 ;
        RECT 50.885 62.855 51.055 63.025 ;
        RECT 51.345 62.855 51.515 63.025 ;
        RECT 51.805 62.855 51.975 63.025 ;
        RECT 52.265 62.855 52.435 63.025 ;
        RECT 52.725 62.855 52.895 63.025 ;
        RECT 53.185 62.855 53.355 63.025 ;
        RECT 53.645 62.855 53.815 63.025 ;
        RECT 54.105 62.855 54.275 63.025 ;
        RECT 54.565 62.855 54.735 63.025 ;
        RECT 55.025 62.855 55.195 63.025 ;
        RECT 55.485 62.855 55.655 63.025 ;
        RECT 55.945 62.855 56.115 63.025 ;
        RECT 56.405 62.855 56.575 63.025 ;
        RECT 56.865 62.855 57.035 63.025 ;
        RECT 57.325 62.855 57.495 63.025 ;
        RECT 57.785 62.855 57.955 63.025 ;
        RECT 58.245 62.855 58.415 63.025 ;
        RECT 58.705 62.855 58.875 63.025 ;
        RECT 59.165 62.855 59.335 63.025 ;
        RECT 59.625 62.855 59.795 63.025 ;
        RECT 60.085 62.855 60.255 63.025 ;
        RECT 60.545 62.855 60.715 63.025 ;
        RECT 61.005 62.855 61.175 63.025 ;
        RECT 61.465 62.855 61.635 63.025 ;
        RECT 61.925 62.855 62.095 63.025 ;
        RECT 62.385 62.855 62.555 63.025 ;
        RECT 62.845 62.855 63.015 63.025 ;
        RECT 63.305 62.855 63.475 63.025 ;
        RECT 63.765 62.855 63.935 63.025 ;
        RECT 64.225 62.855 64.395 63.025 ;
        RECT 64.685 62.855 64.855 63.025 ;
        RECT 65.145 62.855 65.315 63.025 ;
        RECT 65.605 62.855 65.775 63.025 ;
        RECT 66.065 62.855 66.235 63.025 ;
        RECT 66.525 62.855 66.695 63.025 ;
        RECT 66.985 62.855 67.155 63.025 ;
        RECT 67.445 62.855 67.615 63.025 ;
        RECT 67.905 62.855 68.075 63.025 ;
        RECT 68.365 62.855 68.535 63.025 ;
        RECT 68.825 62.855 68.995 63.025 ;
        RECT 69.285 62.855 69.455 63.025 ;
        RECT 69.745 62.855 69.915 63.025 ;
        RECT 70.205 62.855 70.375 63.025 ;
        RECT 70.665 62.855 70.835 63.025 ;
        RECT 71.125 62.855 71.295 63.025 ;
        RECT 71.585 62.855 71.755 63.025 ;
        RECT 72.045 62.855 72.215 63.025 ;
        RECT 72.505 62.855 72.675 63.025 ;
        RECT 72.965 62.855 73.135 63.025 ;
        RECT 73.425 62.855 73.595 63.025 ;
        RECT 73.885 62.855 74.055 63.025 ;
        RECT 74.345 62.855 74.515 63.025 ;
        RECT 74.805 62.855 74.975 63.025 ;
        RECT 75.265 62.855 75.435 63.025 ;
        RECT 75.725 62.855 75.895 63.025 ;
        RECT 76.185 62.855 76.355 63.025 ;
        RECT 76.645 62.855 76.815 63.025 ;
        RECT 77.105 62.855 77.275 63.025 ;
        RECT 77.565 62.855 77.735 63.025 ;
        RECT 78.025 62.855 78.195 63.025 ;
        RECT 78.485 62.855 78.655 63.025 ;
        RECT 78.945 62.855 79.115 63.025 ;
        RECT 79.405 62.855 79.575 63.025 ;
        RECT 79.865 62.855 80.035 63.025 ;
        RECT 80.325 62.855 80.495 63.025 ;
        RECT 80.785 62.855 80.955 63.025 ;
        RECT 81.245 62.855 81.415 63.025 ;
        RECT 81.705 62.855 81.875 63.025 ;
        RECT 82.165 62.855 82.335 63.025 ;
        RECT 82.625 62.855 82.795 63.025 ;
        RECT 83.085 62.855 83.255 63.025 ;
        RECT 83.545 62.855 83.715 63.025 ;
        RECT 84.005 62.855 84.175 63.025 ;
        RECT 84.465 62.855 84.635 63.025 ;
        RECT 84.925 62.855 85.095 63.025 ;
        RECT 85.385 62.855 85.555 63.025 ;
        RECT 85.845 62.855 86.015 63.025 ;
        RECT 86.305 62.855 86.475 63.025 ;
        RECT 86.765 62.855 86.935 63.025 ;
        RECT 87.225 62.855 87.395 63.025 ;
        RECT 87.685 62.855 87.855 63.025 ;
        RECT 88.145 62.855 88.315 63.025 ;
        RECT 88.605 62.855 88.775 63.025 ;
        RECT 89.065 62.855 89.235 63.025 ;
        RECT 89.525 62.855 89.695 63.025 ;
        RECT 89.985 62.855 90.155 63.025 ;
        RECT 90.445 62.855 90.615 63.025 ;
        RECT 90.905 62.855 91.075 63.025 ;
        RECT 91.365 62.855 91.535 63.025 ;
        RECT 91.825 62.855 91.995 63.025 ;
        RECT 92.285 62.855 92.455 63.025 ;
        RECT 92.745 62.855 92.915 63.025 ;
        RECT 93.205 62.855 93.375 63.025 ;
        RECT 93.665 62.855 93.835 63.025 ;
        RECT 94.125 62.855 94.295 63.025 ;
        RECT 94.585 62.855 94.755 63.025 ;
        RECT 95.045 62.855 95.215 63.025 ;
        RECT 95.505 62.855 95.675 63.025 ;
        RECT 95.965 62.855 96.135 63.025 ;
        RECT 96.425 62.855 96.595 63.025 ;
        RECT 96.885 62.855 97.055 63.025 ;
        RECT 97.345 62.855 97.515 63.025 ;
        RECT 97.805 62.855 97.975 63.025 ;
        RECT 98.265 62.855 98.435 63.025 ;
        RECT 98.725 62.855 98.895 63.025 ;
        RECT 99.185 62.855 99.355 63.025 ;
        RECT 99.645 62.855 99.815 63.025 ;
        RECT 16.845 57.415 17.015 57.585 ;
        RECT 17.305 57.415 17.475 57.585 ;
        RECT 17.765 57.415 17.935 57.585 ;
        RECT 18.225 57.415 18.395 57.585 ;
        RECT 18.685 57.415 18.855 57.585 ;
        RECT 19.145 57.415 19.315 57.585 ;
        RECT 19.605 57.415 19.775 57.585 ;
        RECT 20.065 57.415 20.235 57.585 ;
        RECT 20.525 57.415 20.695 57.585 ;
        RECT 20.985 57.415 21.155 57.585 ;
        RECT 21.445 57.415 21.615 57.585 ;
        RECT 21.905 57.415 22.075 57.585 ;
        RECT 22.365 57.415 22.535 57.585 ;
        RECT 22.825 57.415 22.995 57.585 ;
        RECT 23.285 57.415 23.455 57.585 ;
        RECT 23.745 57.415 23.915 57.585 ;
        RECT 24.205 57.415 24.375 57.585 ;
        RECT 24.665 57.415 24.835 57.585 ;
        RECT 25.125 57.415 25.295 57.585 ;
        RECT 25.585 57.415 25.755 57.585 ;
        RECT 26.045 57.415 26.215 57.585 ;
        RECT 26.505 57.415 26.675 57.585 ;
        RECT 26.965 57.415 27.135 57.585 ;
        RECT 27.425 57.415 27.595 57.585 ;
        RECT 27.885 57.415 28.055 57.585 ;
        RECT 28.345 57.415 28.515 57.585 ;
        RECT 28.805 57.415 28.975 57.585 ;
        RECT 29.265 57.415 29.435 57.585 ;
        RECT 29.725 57.415 29.895 57.585 ;
        RECT 30.185 57.415 30.355 57.585 ;
        RECT 30.645 57.415 30.815 57.585 ;
        RECT 31.105 57.415 31.275 57.585 ;
        RECT 31.565 57.415 31.735 57.585 ;
        RECT 32.025 57.415 32.195 57.585 ;
        RECT 32.485 57.415 32.655 57.585 ;
        RECT 32.945 57.415 33.115 57.585 ;
        RECT 33.405 57.415 33.575 57.585 ;
        RECT 33.865 57.415 34.035 57.585 ;
        RECT 34.325 57.415 34.495 57.585 ;
        RECT 34.785 57.415 34.955 57.585 ;
        RECT 35.245 57.415 35.415 57.585 ;
        RECT 35.705 57.415 35.875 57.585 ;
        RECT 36.165 57.415 36.335 57.585 ;
        RECT 36.625 57.415 36.795 57.585 ;
        RECT 37.085 57.415 37.255 57.585 ;
        RECT 37.545 57.415 37.715 57.585 ;
        RECT 38.005 57.415 38.175 57.585 ;
        RECT 38.465 57.415 38.635 57.585 ;
        RECT 38.925 57.415 39.095 57.585 ;
        RECT 39.385 57.415 39.555 57.585 ;
        RECT 39.845 57.415 40.015 57.585 ;
        RECT 40.305 57.415 40.475 57.585 ;
        RECT 40.765 57.415 40.935 57.585 ;
        RECT 41.225 57.415 41.395 57.585 ;
        RECT 41.685 57.415 41.855 57.585 ;
        RECT 42.145 57.415 42.315 57.585 ;
        RECT 42.605 57.415 42.775 57.585 ;
        RECT 43.065 57.415 43.235 57.585 ;
        RECT 43.525 57.415 43.695 57.585 ;
        RECT 43.985 57.415 44.155 57.585 ;
        RECT 44.445 57.415 44.615 57.585 ;
        RECT 44.905 57.415 45.075 57.585 ;
        RECT 45.365 57.415 45.535 57.585 ;
        RECT 45.825 57.415 45.995 57.585 ;
        RECT 46.285 57.415 46.455 57.585 ;
        RECT 46.745 57.415 46.915 57.585 ;
        RECT 47.205 57.415 47.375 57.585 ;
        RECT 47.665 57.415 47.835 57.585 ;
        RECT 48.125 57.415 48.295 57.585 ;
        RECT 48.585 57.415 48.755 57.585 ;
        RECT 49.045 57.415 49.215 57.585 ;
        RECT 49.505 57.415 49.675 57.585 ;
        RECT 49.965 57.415 50.135 57.585 ;
        RECT 50.425 57.415 50.595 57.585 ;
        RECT 50.885 57.415 51.055 57.585 ;
        RECT 51.345 57.415 51.515 57.585 ;
        RECT 51.805 57.415 51.975 57.585 ;
        RECT 52.265 57.415 52.435 57.585 ;
        RECT 52.725 57.415 52.895 57.585 ;
        RECT 53.185 57.415 53.355 57.585 ;
        RECT 53.645 57.415 53.815 57.585 ;
        RECT 54.105 57.415 54.275 57.585 ;
        RECT 54.565 57.415 54.735 57.585 ;
        RECT 55.025 57.415 55.195 57.585 ;
        RECT 55.485 57.415 55.655 57.585 ;
        RECT 55.945 57.415 56.115 57.585 ;
        RECT 56.405 57.415 56.575 57.585 ;
        RECT 56.865 57.415 57.035 57.585 ;
        RECT 57.325 57.415 57.495 57.585 ;
        RECT 57.785 57.415 57.955 57.585 ;
        RECT 58.245 57.415 58.415 57.585 ;
        RECT 58.705 57.415 58.875 57.585 ;
        RECT 59.165 57.415 59.335 57.585 ;
        RECT 59.625 57.415 59.795 57.585 ;
        RECT 60.085 57.415 60.255 57.585 ;
        RECT 60.545 57.415 60.715 57.585 ;
        RECT 61.005 57.415 61.175 57.585 ;
        RECT 61.465 57.415 61.635 57.585 ;
        RECT 61.925 57.415 62.095 57.585 ;
        RECT 62.385 57.415 62.555 57.585 ;
        RECT 62.845 57.415 63.015 57.585 ;
        RECT 63.305 57.415 63.475 57.585 ;
        RECT 63.765 57.415 63.935 57.585 ;
        RECT 64.225 57.415 64.395 57.585 ;
        RECT 64.685 57.415 64.855 57.585 ;
        RECT 65.145 57.415 65.315 57.585 ;
        RECT 65.605 57.415 65.775 57.585 ;
        RECT 66.065 57.415 66.235 57.585 ;
        RECT 66.525 57.415 66.695 57.585 ;
        RECT 66.985 57.415 67.155 57.585 ;
        RECT 67.445 57.415 67.615 57.585 ;
        RECT 67.905 57.415 68.075 57.585 ;
        RECT 68.365 57.415 68.535 57.585 ;
        RECT 68.825 57.415 68.995 57.585 ;
        RECT 69.285 57.415 69.455 57.585 ;
        RECT 69.745 57.415 69.915 57.585 ;
        RECT 70.205 57.415 70.375 57.585 ;
        RECT 70.665 57.415 70.835 57.585 ;
        RECT 71.125 57.415 71.295 57.585 ;
        RECT 71.585 57.415 71.755 57.585 ;
        RECT 72.045 57.415 72.215 57.585 ;
        RECT 72.505 57.415 72.675 57.585 ;
        RECT 72.965 57.415 73.135 57.585 ;
        RECT 73.425 57.415 73.595 57.585 ;
        RECT 73.885 57.415 74.055 57.585 ;
        RECT 74.345 57.415 74.515 57.585 ;
        RECT 74.805 57.415 74.975 57.585 ;
        RECT 75.265 57.415 75.435 57.585 ;
        RECT 75.725 57.415 75.895 57.585 ;
        RECT 76.185 57.415 76.355 57.585 ;
        RECT 76.645 57.415 76.815 57.585 ;
        RECT 77.105 57.415 77.275 57.585 ;
        RECT 77.565 57.415 77.735 57.585 ;
        RECT 78.025 57.415 78.195 57.585 ;
        RECT 78.485 57.415 78.655 57.585 ;
        RECT 78.945 57.415 79.115 57.585 ;
        RECT 79.405 57.415 79.575 57.585 ;
        RECT 79.865 57.415 80.035 57.585 ;
        RECT 80.325 57.415 80.495 57.585 ;
        RECT 80.785 57.415 80.955 57.585 ;
        RECT 81.245 57.415 81.415 57.585 ;
        RECT 81.705 57.415 81.875 57.585 ;
        RECT 82.165 57.415 82.335 57.585 ;
        RECT 82.625 57.415 82.795 57.585 ;
        RECT 83.085 57.415 83.255 57.585 ;
        RECT 83.545 57.415 83.715 57.585 ;
        RECT 84.005 57.415 84.175 57.585 ;
        RECT 84.465 57.415 84.635 57.585 ;
        RECT 84.925 57.415 85.095 57.585 ;
        RECT 85.385 57.415 85.555 57.585 ;
        RECT 85.845 57.415 86.015 57.585 ;
        RECT 86.305 57.415 86.475 57.585 ;
        RECT 86.765 57.415 86.935 57.585 ;
        RECT 87.225 57.415 87.395 57.585 ;
        RECT 87.685 57.415 87.855 57.585 ;
        RECT 88.145 57.415 88.315 57.585 ;
        RECT 88.605 57.415 88.775 57.585 ;
        RECT 89.065 57.415 89.235 57.585 ;
        RECT 89.525 57.415 89.695 57.585 ;
        RECT 89.985 57.415 90.155 57.585 ;
        RECT 90.445 57.415 90.615 57.585 ;
        RECT 90.905 57.415 91.075 57.585 ;
        RECT 91.365 57.415 91.535 57.585 ;
        RECT 91.825 57.415 91.995 57.585 ;
        RECT 92.285 57.415 92.455 57.585 ;
        RECT 92.745 57.415 92.915 57.585 ;
        RECT 93.205 57.415 93.375 57.585 ;
        RECT 93.665 57.415 93.835 57.585 ;
        RECT 94.125 57.415 94.295 57.585 ;
        RECT 94.585 57.415 94.755 57.585 ;
        RECT 95.045 57.415 95.215 57.585 ;
        RECT 95.505 57.415 95.675 57.585 ;
        RECT 95.965 57.415 96.135 57.585 ;
        RECT 96.425 57.415 96.595 57.585 ;
        RECT 96.885 57.415 97.055 57.585 ;
        RECT 97.345 57.415 97.515 57.585 ;
        RECT 97.805 57.415 97.975 57.585 ;
        RECT 98.265 57.415 98.435 57.585 ;
        RECT 98.725 57.415 98.895 57.585 ;
        RECT 99.185 57.415 99.355 57.585 ;
        RECT 99.645 57.415 99.815 57.585 ;
        RECT 16.845 51.975 17.015 52.145 ;
        RECT 17.305 51.975 17.475 52.145 ;
        RECT 17.765 51.975 17.935 52.145 ;
        RECT 18.225 51.975 18.395 52.145 ;
        RECT 18.685 51.975 18.855 52.145 ;
        RECT 19.145 51.975 19.315 52.145 ;
        RECT 19.605 51.975 19.775 52.145 ;
        RECT 20.065 51.975 20.235 52.145 ;
        RECT 20.525 51.975 20.695 52.145 ;
        RECT 20.985 51.975 21.155 52.145 ;
        RECT 21.445 51.975 21.615 52.145 ;
        RECT 21.905 51.975 22.075 52.145 ;
        RECT 22.365 51.975 22.535 52.145 ;
        RECT 22.825 51.975 22.995 52.145 ;
        RECT 23.285 51.975 23.455 52.145 ;
        RECT 23.745 51.975 23.915 52.145 ;
        RECT 24.205 51.975 24.375 52.145 ;
        RECT 24.665 51.975 24.835 52.145 ;
        RECT 25.125 51.975 25.295 52.145 ;
        RECT 25.585 51.975 25.755 52.145 ;
        RECT 26.045 51.975 26.215 52.145 ;
        RECT 26.505 51.975 26.675 52.145 ;
        RECT 26.965 51.975 27.135 52.145 ;
        RECT 27.425 51.975 27.595 52.145 ;
        RECT 27.885 51.975 28.055 52.145 ;
        RECT 28.345 51.975 28.515 52.145 ;
        RECT 28.805 51.975 28.975 52.145 ;
        RECT 29.265 51.975 29.435 52.145 ;
        RECT 29.725 51.975 29.895 52.145 ;
        RECT 30.185 51.975 30.355 52.145 ;
        RECT 30.645 51.975 30.815 52.145 ;
        RECT 31.105 51.975 31.275 52.145 ;
        RECT 31.565 51.975 31.735 52.145 ;
        RECT 32.025 51.975 32.195 52.145 ;
        RECT 32.485 51.975 32.655 52.145 ;
        RECT 32.945 51.975 33.115 52.145 ;
        RECT 33.405 51.975 33.575 52.145 ;
        RECT 33.865 51.975 34.035 52.145 ;
        RECT 34.325 51.975 34.495 52.145 ;
        RECT 34.785 51.975 34.955 52.145 ;
        RECT 35.245 51.975 35.415 52.145 ;
        RECT 35.705 51.975 35.875 52.145 ;
        RECT 36.165 51.975 36.335 52.145 ;
        RECT 36.625 51.975 36.795 52.145 ;
        RECT 37.085 51.975 37.255 52.145 ;
        RECT 37.545 51.975 37.715 52.145 ;
        RECT 38.005 51.975 38.175 52.145 ;
        RECT 38.465 51.975 38.635 52.145 ;
        RECT 38.925 51.975 39.095 52.145 ;
        RECT 39.385 51.975 39.555 52.145 ;
        RECT 39.845 51.975 40.015 52.145 ;
        RECT 40.305 51.975 40.475 52.145 ;
        RECT 40.765 51.975 40.935 52.145 ;
        RECT 41.225 51.975 41.395 52.145 ;
        RECT 41.685 51.975 41.855 52.145 ;
        RECT 42.145 51.975 42.315 52.145 ;
        RECT 42.605 51.975 42.775 52.145 ;
        RECT 43.065 51.975 43.235 52.145 ;
        RECT 43.525 51.975 43.695 52.145 ;
        RECT 43.985 51.975 44.155 52.145 ;
        RECT 44.445 51.975 44.615 52.145 ;
        RECT 44.905 51.975 45.075 52.145 ;
        RECT 45.365 51.975 45.535 52.145 ;
        RECT 45.825 51.975 45.995 52.145 ;
        RECT 46.285 51.975 46.455 52.145 ;
        RECT 46.745 51.975 46.915 52.145 ;
        RECT 47.205 51.975 47.375 52.145 ;
        RECT 47.665 51.975 47.835 52.145 ;
        RECT 48.125 51.975 48.295 52.145 ;
        RECT 48.585 51.975 48.755 52.145 ;
        RECT 49.045 51.975 49.215 52.145 ;
        RECT 49.505 51.975 49.675 52.145 ;
        RECT 49.965 51.975 50.135 52.145 ;
        RECT 50.425 51.975 50.595 52.145 ;
        RECT 50.885 51.975 51.055 52.145 ;
        RECT 51.345 51.975 51.515 52.145 ;
        RECT 51.805 51.975 51.975 52.145 ;
        RECT 52.265 51.975 52.435 52.145 ;
        RECT 52.725 51.975 52.895 52.145 ;
        RECT 53.185 51.975 53.355 52.145 ;
        RECT 53.645 51.975 53.815 52.145 ;
        RECT 54.105 51.975 54.275 52.145 ;
        RECT 54.565 51.975 54.735 52.145 ;
        RECT 55.025 51.975 55.195 52.145 ;
        RECT 55.485 51.975 55.655 52.145 ;
        RECT 55.945 51.975 56.115 52.145 ;
        RECT 56.405 51.975 56.575 52.145 ;
        RECT 56.865 51.975 57.035 52.145 ;
        RECT 57.325 51.975 57.495 52.145 ;
        RECT 57.785 51.975 57.955 52.145 ;
        RECT 58.245 51.975 58.415 52.145 ;
        RECT 58.705 51.975 58.875 52.145 ;
        RECT 59.165 51.975 59.335 52.145 ;
        RECT 59.625 51.975 59.795 52.145 ;
        RECT 60.085 51.975 60.255 52.145 ;
        RECT 60.545 51.975 60.715 52.145 ;
        RECT 61.005 51.975 61.175 52.145 ;
        RECT 61.465 51.975 61.635 52.145 ;
        RECT 61.925 51.975 62.095 52.145 ;
        RECT 62.385 51.975 62.555 52.145 ;
        RECT 62.845 51.975 63.015 52.145 ;
        RECT 63.305 51.975 63.475 52.145 ;
        RECT 63.765 51.975 63.935 52.145 ;
        RECT 64.225 51.975 64.395 52.145 ;
        RECT 64.685 51.975 64.855 52.145 ;
        RECT 65.145 51.975 65.315 52.145 ;
        RECT 65.605 51.975 65.775 52.145 ;
        RECT 66.065 51.975 66.235 52.145 ;
        RECT 66.525 51.975 66.695 52.145 ;
        RECT 66.985 51.975 67.155 52.145 ;
        RECT 67.445 51.975 67.615 52.145 ;
        RECT 67.905 51.975 68.075 52.145 ;
        RECT 68.365 51.975 68.535 52.145 ;
        RECT 68.825 51.975 68.995 52.145 ;
        RECT 69.285 51.975 69.455 52.145 ;
        RECT 69.745 51.975 69.915 52.145 ;
        RECT 70.205 51.975 70.375 52.145 ;
        RECT 70.665 51.975 70.835 52.145 ;
        RECT 71.125 51.975 71.295 52.145 ;
        RECT 71.585 51.975 71.755 52.145 ;
        RECT 72.045 51.975 72.215 52.145 ;
        RECT 72.505 51.975 72.675 52.145 ;
        RECT 72.965 51.975 73.135 52.145 ;
        RECT 73.425 51.975 73.595 52.145 ;
        RECT 73.885 51.975 74.055 52.145 ;
        RECT 74.345 51.975 74.515 52.145 ;
        RECT 74.805 51.975 74.975 52.145 ;
        RECT 75.265 51.975 75.435 52.145 ;
        RECT 75.725 51.975 75.895 52.145 ;
        RECT 76.185 51.975 76.355 52.145 ;
        RECT 76.645 51.975 76.815 52.145 ;
        RECT 77.105 51.975 77.275 52.145 ;
        RECT 77.565 51.975 77.735 52.145 ;
        RECT 78.025 51.975 78.195 52.145 ;
        RECT 78.485 51.975 78.655 52.145 ;
        RECT 78.945 51.975 79.115 52.145 ;
        RECT 79.405 51.975 79.575 52.145 ;
        RECT 79.865 51.975 80.035 52.145 ;
        RECT 80.325 51.975 80.495 52.145 ;
        RECT 80.785 51.975 80.955 52.145 ;
        RECT 81.245 51.975 81.415 52.145 ;
        RECT 81.705 51.975 81.875 52.145 ;
        RECT 82.165 51.975 82.335 52.145 ;
        RECT 82.625 51.975 82.795 52.145 ;
        RECT 83.085 51.975 83.255 52.145 ;
        RECT 83.545 51.975 83.715 52.145 ;
        RECT 84.005 51.975 84.175 52.145 ;
        RECT 84.465 51.975 84.635 52.145 ;
        RECT 84.925 51.975 85.095 52.145 ;
        RECT 85.385 51.975 85.555 52.145 ;
        RECT 85.845 51.975 86.015 52.145 ;
        RECT 86.305 51.975 86.475 52.145 ;
        RECT 86.765 51.975 86.935 52.145 ;
        RECT 87.225 51.975 87.395 52.145 ;
        RECT 87.685 51.975 87.855 52.145 ;
        RECT 88.145 51.975 88.315 52.145 ;
        RECT 88.605 51.975 88.775 52.145 ;
        RECT 89.065 51.975 89.235 52.145 ;
        RECT 89.525 51.975 89.695 52.145 ;
        RECT 89.985 51.975 90.155 52.145 ;
        RECT 90.445 51.975 90.615 52.145 ;
        RECT 90.905 51.975 91.075 52.145 ;
        RECT 91.365 51.975 91.535 52.145 ;
        RECT 91.825 51.975 91.995 52.145 ;
        RECT 92.285 51.975 92.455 52.145 ;
        RECT 92.745 51.975 92.915 52.145 ;
        RECT 93.205 51.975 93.375 52.145 ;
        RECT 93.665 51.975 93.835 52.145 ;
        RECT 94.125 51.975 94.295 52.145 ;
        RECT 94.585 51.975 94.755 52.145 ;
        RECT 95.045 51.975 95.215 52.145 ;
        RECT 95.505 51.975 95.675 52.145 ;
        RECT 95.965 51.975 96.135 52.145 ;
        RECT 96.425 51.975 96.595 52.145 ;
        RECT 96.885 51.975 97.055 52.145 ;
        RECT 97.345 51.975 97.515 52.145 ;
        RECT 97.805 51.975 97.975 52.145 ;
        RECT 98.265 51.975 98.435 52.145 ;
        RECT 98.725 51.975 98.895 52.145 ;
        RECT 99.185 51.975 99.355 52.145 ;
        RECT 99.645 51.975 99.815 52.145 ;
        RECT 16.845 46.535 17.015 46.705 ;
        RECT 17.305 46.535 17.475 46.705 ;
        RECT 17.765 46.535 17.935 46.705 ;
        RECT 18.225 46.535 18.395 46.705 ;
        RECT 18.685 46.535 18.855 46.705 ;
        RECT 19.145 46.535 19.315 46.705 ;
        RECT 19.605 46.535 19.775 46.705 ;
        RECT 20.065 46.535 20.235 46.705 ;
        RECT 20.525 46.535 20.695 46.705 ;
        RECT 20.985 46.535 21.155 46.705 ;
        RECT 21.445 46.535 21.615 46.705 ;
        RECT 21.905 46.535 22.075 46.705 ;
        RECT 22.365 46.535 22.535 46.705 ;
        RECT 22.825 46.535 22.995 46.705 ;
        RECT 23.285 46.535 23.455 46.705 ;
        RECT 23.745 46.535 23.915 46.705 ;
        RECT 24.205 46.535 24.375 46.705 ;
        RECT 24.665 46.535 24.835 46.705 ;
        RECT 25.125 46.535 25.295 46.705 ;
        RECT 25.585 46.535 25.755 46.705 ;
        RECT 26.045 46.535 26.215 46.705 ;
        RECT 26.505 46.535 26.675 46.705 ;
        RECT 26.965 46.535 27.135 46.705 ;
        RECT 27.425 46.535 27.595 46.705 ;
        RECT 27.885 46.535 28.055 46.705 ;
        RECT 28.345 46.535 28.515 46.705 ;
        RECT 28.805 46.535 28.975 46.705 ;
        RECT 29.265 46.535 29.435 46.705 ;
        RECT 29.725 46.535 29.895 46.705 ;
        RECT 30.185 46.535 30.355 46.705 ;
        RECT 30.645 46.535 30.815 46.705 ;
        RECT 31.105 46.535 31.275 46.705 ;
        RECT 31.565 46.535 31.735 46.705 ;
        RECT 32.025 46.535 32.195 46.705 ;
        RECT 32.485 46.535 32.655 46.705 ;
        RECT 32.945 46.535 33.115 46.705 ;
        RECT 33.405 46.535 33.575 46.705 ;
        RECT 33.865 46.535 34.035 46.705 ;
        RECT 34.325 46.535 34.495 46.705 ;
        RECT 34.785 46.535 34.955 46.705 ;
        RECT 35.245 46.535 35.415 46.705 ;
        RECT 35.705 46.535 35.875 46.705 ;
        RECT 36.165 46.535 36.335 46.705 ;
        RECT 36.625 46.535 36.795 46.705 ;
        RECT 37.085 46.535 37.255 46.705 ;
        RECT 37.545 46.535 37.715 46.705 ;
        RECT 38.005 46.535 38.175 46.705 ;
        RECT 38.465 46.535 38.635 46.705 ;
        RECT 38.925 46.535 39.095 46.705 ;
        RECT 39.385 46.535 39.555 46.705 ;
        RECT 39.845 46.535 40.015 46.705 ;
        RECT 40.305 46.535 40.475 46.705 ;
        RECT 40.765 46.535 40.935 46.705 ;
        RECT 41.225 46.535 41.395 46.705 ;
        RECT 41.685 46.535 41.855 46.705 ;
        RECT 42.145 46.535 42.315 46.705 ;
        RECT 42.605 46.535 42.775 46.705 ;
        RECT 43.065 46.535 43.235 46.705 ;
        RECT 43.525 46.535 43.695 46.705 ;
        RECT 43.985 46.535 44.155 46.705 ;
        RECT 44.445 46.535 44.615 46.705 ;
        RECT 44.905 46.535 45.075 46.705 ;
        RECT 45.365 46.535 45.535 46.705 ;
        RECT 45.825 46.535 45.995 46.705 ;
        RECT 46.285 46.535 46.455 46.705 ;
        RECT 46.745 46.535 46.915 46.705 ;
        RECT 47.205 46.535 47.375 46.705 ;
        RECT 47.665 46.535 47.835 46.705 ;
        RECT 48.125 46.535 48.295 46.705 ;
        RECT 48.585 46.535 48.755 46.705 ;
        RECT 49.045 46.535 49.215 46.705 ;
        RECT 49.505 46.535 49.675 46.705 ;
        RECT 49.965 46.535 50.135 46.705 ;
        RECT 50.425 46.535 50.595 46.705 ;
        RECT 50.885 46.535 51.055 46.705 ;
        RECT 51.345 46.535 51.515 46.705 ;
        RECT 51.805 46.535 51.975 46.705 ;
        RECT 52.265 46.535 52.435 46.705 ;
        RECT 52.725 46.535 52.895 46.705 ;
        RECT 53.185 46.535 53.355 46.705 ;
        RECT 53.645 46.535 53.815 46.705 ;
        RECT 54.105 46.535 54.275 46.705 ;
        RECT 54.565 46.535 54.735 46.705 ;
        RECT 55.025 46.535 55.195 46.705 ;
        RECT 55.485 46.535 55.655 46.705 ;
        RECT 55.945 46.535 56.115 46.705 ;
        RECT 56.405 46.535 56.575 46.705 ;
        RECT 56.865 46.535 57.035 46.705 ;
        RECT 57.325 46.535 57.495 46.705 ;
        RECT 57.785 46.535 57.955 46.705 ;
        RECT 58.245 46.535 58.415 46.705 ;
        RECT 58.705 46.535 58.875 46.705 ;
        RECT 59.165 46.535 59.335 46.705 ;
        RECT 59.625 46.535 59.795 46.705 ;
        RECT 60.085 46.535 60.255 46.705 ;
        RECT 60.545 46.535 60.715 46.705 ;
        RECT 61.005 46.535 61.175 46.705 ;
        RECT 61.465 46.535 61.635 46.705 ;
        RECT 61.925 46.535 62.095 46.705 ;
        RECT 62.385 46.535 62.555 46.705 ;
        RECT 62.845 46.535 63.015 46.705 ;
        RECT 63.305 46.535 63.475 46.705 ;
        RECT 63.765 46.535 63.935 46.705 ;
        RECT 64.225 46.535 64.395 46.705 ;
        RECT 64.685 46.535 64.855 46.705 ;
        RECT 65.145 46.535 65.315 46.705 ;
        RECT 65.605 46.535 65.775 46.705 ;
        RECT 66.065 46.535 66.235 46.705 ;
        RECT 66.525 46.535 66.695 46.705 ;
        RECT 66.985 46.535 67.155 46.705 ;
        RECT 67.445 46.535 67.615 46.705 ;
        RECT 67.905 46.535 68.075 46.705 ;
        RECT 68.365 46.535 68.535 46.705 ;
        RECT 68.825 46.535 68.995 46.705 ;
        RECT 69.285 46.535 69.455 46.705 ;
        RECT 69.745 46.535 69.915 46.705 ;
        RECT 70.205 46.535 70.375 46.705 ;
        RECT 70.665 46.535 70.835 46.705 ;
        RECT 71.125 46.535 71.295 46.705 ;
        RECT 71.585 46.535 71.755 46.705 ;
        RECT 72.045 46.535 72.215 46.705 ;
        RECT 72.505 46.535 72.675 46.705 ;
        RECT 72.965 46.535 73.135 46.705 ;
        RECT 73.425 46.535 73.595 46.705 ;
        RECT 73.885 46.535 74.055 46.705 ;
        RECT 74.345 46.535 74.515 46.705 ;
        RECT 74.805 46.535 74.975 46.705 ;
        RECT 75.265 46.535 75.435 46.705 ;
        RECT 75.725 46.535 75.895 46.705 ;
        RECT 76.185 46.535 76.355 46.705 ;
        RECT 76.645 46.535 76.815 46.705 ;
        RECT 77.105 46.535 77.275 46.705 ;
        RECT 77.565 46.535 77.735 46.705 ;
        RECT 78.025 46.535 78.195 46.705 ;
        RECT 78.485 46.535 78.655 46.705 ;
        RECT 78.945 46.535 79.115 46.705 ;
        RECT 79.405 46.535 79.575 46.705 ;
        RECT 79.865 46.535 80.035 46.705 ;
        RECT 80.325 46.535 80.495 46.705 ;
        RECT 80.785 46.535 80.955 46.705 ;
        RECT 81.245 46.535 81.415 46.705 ;
        RECT 81.705 46.535 81.875 46.705 ;
        RECT 82.165 46.535 82.335 46.705 ;
        RECT 82.625 46.535 82.795 46.705 ;
        RECT 83.085 46.535 83.255 46.705 ;
        RECT 83.545 46.535 83.715 46.705 ;
        RECT 84.005 46.535 84.175 46.705 ;
        RECT 84.465 46.535 84.635 46.705 ;
        RECT 84.925 46.535 85.095 46.705 ;
        RECT 85.385 46.535 85.555 46.705 ;
        RECT 85.845 46.535 86.015 46.705 ;
        RECT 86.305 46.535 86.475 46.705 ;
        RECT 86.765 46.535 86.935 46.705 ;
        RECT 87.225 46.535 87.395 46.705 ;
        RECT 87.685 46.535 87.855 46.705 ;
        RECT 88.145 46.535 88.315 46.705 ;
        RECT 88.605 46.535 88.775 46.705 ;
        RECT 89.065 46.535 89.235 46.705 ;
        RECT 89.525 46.535 89.695 46.705 ;
        RECT 89.985 46.535 90.155 46.705 ;
        RECT 90.445 46.535 90.615 46.705 ;
        RECT 90.905 46.535 91.075 46.705 ;
        RECT 91.365 46.535 91.535 46.705 ;
        RECT 91.825 46.535 91.995 46.705 ;
        RECT 92.285 46.535 92.455 46.705 ;
        RECT 92.745 46.535 92.915 46.705 ;
        RECT 93.205 46.535 93.375 46.705 ;
        RECT 93.665 46.535 93.835 46.705 ;
        RECT 94.125 46.535 94.295 46.705 ;
        RECT 94.585 46.535 94.755 46.705 ;
        RECT 95.045 46.535 95.215 46.705 ;
        RECT 95.505 46.535 95.675 46.705 ;
        RECT 95.965 46.535 96.135 46.705 ;
        RECT 96.425 46.535 96.595 46.705 ;
        RECT 96.885 46.535 97.055 46.705 ;
        RECT 97.345 46.535 97.515 46.705 ;
        RECT 97.805 46.535 97.975 46.705 ;
        RECT 98.265 46.535 98.435 46.705 ;
        RECT 98.725 46.535 98.895 46.705 ;
        RECT 99.185 46.535 99.355 46.705 ;
        RECT 99.645 46.535 99.815 46.705 ;
        RECT 16.845 41.095 17.015 41.265 ;
        RECT 17.305 41.095 17.475 41.265 ;
        RECT 17.765 41.095 17.935 41.265 ;
        RECT 18.225 41.095 18.395 41.265 ;
        RECT 18.685 41.095 18.855 41.265 ;
        RECT 19.145 41.095 19.315 41.265 ;
        RECT 19.605 41.095 19.775 41.265 ;
        RECT 20.065 41.095 20.235 41.265 ;
        RECT 20.525 41.095 20.695 41.265 ;
        RECT 20.985 41.095 21.155 41.265 ;
        RECT 21.445 41.095 21.615 41.265 ;
        RECT 21.905 41.095 22.075 41.265 ;
        RECT 22.365 41.095 22.535 41.265 ;
        RECT 22.825 41.095 22.995 41.265 ;
        RECT 23.285 41.095 23.455 41.265 ;
        RECT 23.745 41.095 23.915 41.265 ;
        RECT 24.205 41.095 24.375 41.265 ;
        RECT 24.665 41.095 24.835 41.265 ;
        RECT 25.125 41.095 25.295 41.265 ;
        RECT 25.585 41.095 25.755 41.265 ;
        RECT 26.045 41.095 26.215 41.265 ;
        RECT 26.505 41.095 26.675 41.265 ;
        RECT 26.965 41.095 27.135 41.265 ;
        RECT 27.425 41.095 27.595 41.265 ;
        RECT 27.885 41.095 28.055 41.265 ;
        RECT 28.345 41.095 28.515 41.265 ;
        RECT 28.805 41.095 28.975 41.265 ;
        RECT 29.265 41.095 29.435 41.265 ;
        RECT 29.725 41.095 29.895 41.265 ;
        RECT 30.185 41.095 30.355 41.265 ;
        RECT 30.645 41.095 30.815 41.265 ;
        RECT 31.105 41.095 31.275 41.265 ;
        RECT 31.565 41.095 31.735 41.265 ;
        RECT 32.025 41.095 32.195 41.265 ;
        RECT 32.485 41.095 32.655 41.265 ;
        RECT 32.945 41.095 33.115 41.265 ;
        RECT 33.405 41.095 33.575 41.265 ;
        RECT 33.865 41.095 34.035 41.265 ;
        RECT 34.325 41.095 34.495 41.265 ;
        RECT 34.785 41.095 34.955 41.265 ;
        RECT 35.245 41.095 35.415 41.265 ;
        RECT 35.705 41.095 35.875 41.265 ;
        RECT 36.165 41.095 36.335 41.265 ;
        RECT 36.625 41.095 36.795 41.265 ;
        RECT 37.085 41.095 37.255 41.265 ;
        RECT 37.545 41.095 37.715 41.265 ;
        RECT 38.005 41.095 38.175 41.265 ;
        RECT 38.465 41.095 38.635 41.265 ;
        RECT 38.925 41.095 39.095 41.265 ;
        RECT 39.385 41.095 39.555 41.265 ;
        RECT 39.845 41.095 40.015 41.265 ;
        RECT 40.305 41.095 40.475 41.265 ;
        RECT 40.765 41.095 40.935 41.265 ;
        RECT 41.225 41.095 41.395 41.265 ;
        RECT 41.685 41.095 41.855 41.265 ;
        RECT 42.145 41.095 42.315 41.265 ;
        RECT 42.605 41.095 42.775 41.265 ;
        RECT 43.065 41.095 43.235 41.265 ;
        RECT 43.525 41.095 43.695 41.265 ;
        RECT 43.985 41.095 44.155 41.265 ;
        RECT 44.445 41.095 44.615 41.265 ;
        RECT 44.905 41.095 45.075 41.265 ;
        RECT 45.365 41.095 45.535 41.265 ;
        RECT 45.825 41.095 45.995 41.265 ;
        RECT 46.285 41.095 46.455 41.265 ;
        RECT 46.745 41.095 46.915 41.265 ;
        RECT 47.205 41.095 47.375 41.265 ;
        RECT 47.665 41.095 47.835 41.265 ;
        RECT 48.125 41.095 48.295 41.265 ;
        RECT 48.585 41.095 48.755 41.265 ;
        RECT 49.045 41.095 49.215 41.265 ;
        RECT 49.505 41.095 49.675 41.265 ;
        RECT 49.965 41.095 50.135 41.265 ;
        RECT 50.425 41.095 50.595 41.265 ;
        RECT 50.885 41.095 51.055 41.265 ;
        RECT 51.345 41.095 51.515 41.265 ;
        RECT 51.805 41.095 51.975 41.265 ;
        RECT 52.265 41.095 52.435 41.265 ;
        RECT 52.725 41.095 52.895 41.265 ;
        RECT 53.185 41.095 53.355 41.265 ;
        RECT 53.645 41.095 53.815 41.265 ;
        RECT 54.105 41.095 54.275 41.265 ;
        RECT 54.565 41.095 54.735 41.265 ;
        RECT 55.025 41.095 55.195 41.265 ;
        RECT 55.485 41.095 55.655 41.265 ;
        RECT 55.945 41.095 56.115 41.265 ;
        RECT 56.405 41.095 56.575 41.265 ;
        RECT 56.865 41.095 57.035 41.265 ;
        RECT 57.325 41.095 57.495 41.265 ;
        RECT 57.785 41.095 57.955 41.265 ;
        RECT 58.245 41.095 58.415 41.265 ;
        RECT 58.705 41.095 58.875 41.265 ;
        RECT 59.165 41.095 59.335 41.265 ;
        RECT 59.625 41.095 59.795 41.265 ;
        RECT 60.085 41.095 60.255 41.265 ;
        RECT 60.545 41.095 60.715 41.265 ;
        RECT 61.005 41.095 61.175 41.265 ;
        RECT 61.465 41.095 61.635 41.265 ;
        RECT 61.925 41.095 62.095 41.265 ;
        RECT 62.385 41.095 62.555 41.265 ;
        RECT 62.845 41.095 63.015 41.265 ;
        RECT 63.305 41.095 63.475 41.265 ;
        RECT 63.765 41.095 63.935 41.265 ;
        RECT 64.225 41.095 64.395 41.265 ;
        RECT 64.685 41.095 64.855 41.265 ;
        RECT 65.145 41.095 65.315 41.265 ;
        RECT 65.605 41.095 65.775 41.265 ;
        RECT 66.065 41.095 66.235 41.265 ;
        RECT 66.525 41.095 66.695 41.265 ;
        RECT 66.985 41.095 67.155 41.265 ;
        RECT 67.445 41.095 67.615 41.265 ;
        RECT 67.905 41.095 68.075 41.265 ;
        RECT 68.365 41.095 68.535 41.265 ;
        RECT 68.825 41.095 68.995 41.265 ;
        RECT 69.285 41.095 69.455 41.265 ;
        RECT 69.745 41.095 69.915 41.265 ;
        RECT 70.205 41.095 70.375 41.265 ;
        RECT 70.665 41.095 70.835 41.265 ;
        RECT 71.125 41.095 71.295 41.265 ;
        RECT 71.585 41.095 71.755 41.265 ;
        RECT 72.045 41.095 72.215 41.265 ;
        RECT 72.505 41.095 72.675 41.265 ;
        RECT 72.965 41.095 73.135 41.265 ;
        RECT 73.425 41.095 73.595 41.265 ;
        RECT 73.885 41.095 74.055 41.265 ;
        RECT 74.345 41.095 74.515 41.265 ;
        RECT 74.805 41.095 74.975 41.265 ;
        RECT 75.265 41.095 75.435 41.265 ;
        RECT 75.725 41.095 75.895 41.265 ;
        RECT 76.185 41.095 76.355 41.265 ;
        RECT 76.645 41.095 76.815 41.265 ;
        RECT 77.105 41.095 77.275 41.265 ;
        RECT 77.565 41.095 77.735 41.265 ;
        RECT 78.025 41.095 78.195 41.265 ;
        RECT 78.485 41.095 78.655 41.265 ;
        RECT 78.945 41.095 79.115 41.265 ;
        RECT 79.405 41.095 79.575 41.265 ;
        RECT 79.865 41.095 80.035 41.265 ;
        RECT 80.325 41.095 80.495 41.265 ;
        RECT 80.785 41.095 80.955 41.265 ;
        RECT 81.245 41.095 81.415 41.265 ;
        RECT 81.705 41.095 81.875 41.265 ;
        RECT 82.165 41.095 82.335 41.265 ;
        RECT 82.625 41.095 82.795 41.265 ;
        RECT 83.085 41.095 83.255 41.265 ;
        RECT 83.545 41.095 83.715 41.265 ;
        RECT 84.005 41.095 84.175 41.265 ;
        RECT 84.465 41.095 84.635 41.265 ;
        RECT 84.925 41.095 85.095 41.265 ;
        RECT 85.385 41.095 85.555 41.265 ;
        RECT 85.845 41.095 86.015 41.265 ;
        RECT 86.305 41.095 86.475 41.265 ;
        RECT 86.765 41.095 86.935 41.265 ;
        RECT 87.225 41.095 87.395 41.265 ;
        RECT 87.685 41.095 87.855 41.265 ;
        RECT 88.145 41.095 88.315 41.265 ;
        RECT 88.605 41.095 88.775 41.265 ;
        RECT 89.065 41.095 89.235 41.265 ;
        RECT 89.525 41.095 89.695 41.265 ;
        RECT 89.985 41.095 90.155 41.265 ;
        RECT 90.445 41.095 90.615 41.265 ;
        RECT 90.905 41.095 91.075 41.265 ;
        RECT 91.365 41.095 91.535 41.265 ;
        RECT 91.825 41.095 91.995 41.265 ;
        RECT 92.285 41.095 92.455 41.265 ;
        RECT 92.745 41.095 92.915 41.265 ;
        RECT 93.205 41.095 93.375 41.265 ;
        RECT 93.665 41.095 93.835 41.265 ;
        RECT 94.125 41.095 94.295 41.265 ;
        RECT 94.585 41.095 94.755 41.265 ;
        RECT 95.045 41.095 95.215 41.265 ;
        RECT 95.505 41.095 95.675 41.265 ;
        RECT 95.965 41.095 96.135 41.265 ;
        RECT 96.425 41.095 96.595 41.265 ;
        RECT 96.885 41.095 97.055 41.265 ;
        RECT 97.345 41.095 97.515 41.265 ;
        RECT 97.805 41.095 97.975 41.265 ;
        RECT 98.265 41.095 98.435 41.265 ;
        RECT 98.725 41.095 98.895 41.265 ;
        RECT 99.185 41.095 99.355 41.265 ;
        RECT 99.645 41.095 99.815 41.265 ;
        RECT 16.845 35.655 17.015 35.825 ;
        RECT 17.305 35.655 17.475 35.825 ;
        RECT 17.765 35.655 17.935 35.825 ;
        RECT 18.225 35.655 18.395 35.825 ;
        RECT 18.685 35.655 18.855 35.825 ;
        RECT 19.145 35.655 19.315 35.825 ;
        RECT 19.605 35.655 19.775 35.825 ;
        RECT 20.065 35.655 20.235 35.825 ;
        RECT 20.525 35.655 20.695 35.825 ;
        RECT 20.985 35.655 21.155 35.825 ;
        RECT 21.445 35.655 21.615 35.825 ;
        RECT 21.905 35.655 22.075 35.825 ;
        RECT 22.365 35.655 22.535 35.825 ;
        RECT 22.825 35.655 22.995 35.825 ;
        RECT 23.285 35.655 23.455 35.825 ;
        RECT 23.745 35.655 23.915 35.825 ;
        RECT 24.205 35.655 24.375 35.825 ;
        RECT 24.665 35.655 24.835 35.825 ;
        RECT 25.125 35.655 25.295 35.825 ;
        RECT 25.585 35.655 25.755 35.825 ;
        RECT 26.045 35.655 26.215 35.825 ;
        RECT 26.505 35.655 26.675 35.825 ;
        RECT 26.965 35.655 27.135 35.825 ;
        RECT 27.425 35.655 27.595 35.825 ;
        RECT 27.885 35.655 28.055 35.825 ;
        RECT 28.345 35.655 28.515 35.825 ;
        RECT 28.805 35.655 28.975 35.825 ;
        RECT 29.265 35.655 29.435 35.825 ;
        RECT 29.725 35.655 29.895 35.825 ;
        RECT 30.185 35.655 30.355 35.825 ;
        RECT 30.645 35.655 30.815 35.825 ;
        RECT 31.105 35.655 31.275 35.825 ;
        RECT 31.565 35.655 31.735 35.825 ;
        RECT 32.025 35.655 32.195 35.825 ;
        RECT 32.485 35.655 32.655 35.825 ;
        RECT 32.945 35.655 33.115 35.825 ;
        RECT 33.405 35.655 33.575 35.825 ;
        RECT 33.865 35.655 34.035 35.825 ;
        RECT 34.325 35.655 34.495 35.825 ;
        RECT 34.785 35.655 34.955 35.825 ;
        RECT 35.245 35.655 35.415 35.825 ;
        RECT 35.705 35.655 35.875 35.825 ;
        RECT 36.165 35.655 36.335 35.825 ;
        RECT 36.625 35.655 36.795 35.825 ;
        RECT 37.085 35.655 37.255 35.825 ;
        RECT 37.545 35.655 37.715 35.825 ;
        RECT 38.005 35.655 38.175 35.825 ;
        RECT 38.465 35.655 38.635 35.825 ;
        RECT 38.925 35.655 39.095 35.825 ;
        RECT 39.385 35.655 39.555 35.825 ;
        RECT 39.845 35.655 40.015 35.825 ;
        RECT 40.305 35.655 40.475 35.825 ;
        RECT 40.765 35.655 40.935 35.825 ;
        RECT 41.225 35.655 41.395 35.825 ;
        RECT 41.685 35.655 41.855 35.825 ;
        RECT 42.145 35.655 42.315 35.825 ;
        RECT 42.605 35.655 42.775 35.825 ;
        RECT 43.065 35.655 43.235 35.825 ;
        RECT 43.525 35.655 43.695 35.825 ;
        RECT 43.985 35.655 44.155 35.825 ;
        RECT 44.445 35.655 44.615 35.825 ;
        RECT 44.905 35.655 45.075 35.825 ;
        RECT 45.365 35.655 45.535 35.825 ;
        RECT 45.825 35.655 45.995 35.825 ;
        RECT 46.285 35.655 46.455 35.825 ;
        RECT 46.745 35.655 46.915 35.825 ;
        RECT 47.205 35.655 47.375 35.825 ;
        RECT 47.665 35.655 47.835 35.825 ;
        RECT 48.125 35.655 48.295 35.825 ;
        RECT 48.585 35.655 48.755 35.825 ;
        RECT 49.045 35.655 49.215 35.825 ;
        RECT 49.505 35.655 49.675 35.825 ;
        RECT 49.965 35.655 50.135 35.825 ;
        RECT 50.425 35.655 50.595 35.825 ;
        RECT 50.885 35.655 51.055 35.825 ;
        RECT 51.345 35.655 51.515 35.825 ;
        RECT 51.805 35.655 51.975 35.825 ;
        RECT 52.265 35.655 52.435 35.825 ;
        RECT 52.725 35.655 52.895 35.825 ;
        RECT 53.185 35.655 53.355 35.825 ;
        RECT 53.645 35.655 53.815 35.825 ;
        RECT 54.105 35.655 54.275 35.825 ;
        RECT 54.565 35.655 54.735 35.825 ;
        RECT 55.025 35.655 55.195 35.825 ;
        RECT 55.485 35.655 55.655 35.825 ;
        RECT 55.945 35.655 56.115 35.825 ;
        RECT 56.405 35.655 56.575 35.825 ;
        RECT 56.865 35.655 57.035 35.825 ;
        RECT 57.325 35.655 57.495 35.825 ;
        RECT 57.785 35.655 57.955 35.825 ;
        RECT 58.245 35.655 58.415 35.825 ;
        RECT 58.705 35.655 58.875 35.825 ;
        RECT 59.165 35.655 59.335 35.825 ;
        RECT 59.625 35.655 59.795 35.825 ;
        RECT 60.085 35.655 60.255 35.825 ;
        RECT 60.545 35.655 60.715 35.825 ;
        RECT 61.005 35.655 61.175 35.825 ;
        RECT 61.465 35.655 61.635 35.825 ;
        RECT 61.925 35.655 62.095 35.825 ;
        RECT 62.385 35.655 62.555 35.825 ;
        RECT 62.845 35.655 63.015 35.825 ;
        RECT 63.305 35.655 63.475 35.825 ;
        RECT 63.765 35.655 63.935 35.825 ;
        RECT 64.225 35.655 64.395 35.825 ;
        RECT 64.685 35.655 64.855 35.825 ;
        RECT 65.145 35.655 65.315 35.825 ;
        RECT 65.605 35.655 65.775 35.825 ;
        RECT 66.065 35.655 66.235 35.825 ;
        RECT 66.525 35.655 66.695 35.825 ;
        RECT 66.985 35.655 67.155 35.825 ;
        RECT 67.445 35.655 67.615 35.825 ;
        RECT 67.905 35.655 68.075 35.825 ;
        RECT 68.365 35.655 68.535 35.825 ;
        RECT 68.825 35.655 68.995 35.825 ;
        RECT 69.285 35.655 69.455 35.825 ;
        RECT 69.745 35.655 69.915 35.825 ;
        RECT 70.205 35.655 70.375 35.825 ;
        RECT 70.665 35.655 70.835 35.825 ;
        RECT 71.125 35.655 71.295 35.825 ;
        RECT 71.585 35.655 71.755 35.825 ;
        RECT 72.045 35.655 72.215 35.825 ;
        RECT 72.505 35.655 72.675 35.825 ;
        RECT 72.965 35.655 73.135 35.825 ;
        RECT 73.425 35.655 73.595 35.825 ;
        RECT 73.885 35.655 74.055 35.825 ;
        RECT 74.345 35.655 74.515 35.825 ;
        RECT 74.805 35.655 74.975 35.825 ;
        RECT 75.265 35.655 75.435 35.825 ;
        RECT 75.725 35.655 75.895 35.825 ;
        RECT 76.185 35.655 76.355 35.825 ;
        RECT 76.645 35.655 76.815 35.825 ;
        RECT 77.105 35.655 77.275 35.825 ;
        RECT 77.565 35.655 77.735 35.825 ;
        RECT 78.025 35.655 78.195 35.825 ;
        RECT 78.485 35.655 78.655 35.825 ;
        RECT 78.945 35.655 79.115 35.825 ;
        RECT 79.405 35.655 79.575 35.825 ;
        RECT 79.865 35.655 80.035 35.825 ;
        RECT 80.325 35.655 80.495 35.825 ;
        RECT 80.785 35.655 80.955 35.825 ;
        RECT 81.245 35.655 81.415 35.825 ;
        RECT 81.705 35.655 81.875 35.825 ;
        RECT 82.165 35.655 82.335 35.825 ;
        RECT 82.625 35.655 82.795 35.825 ;
        RECT 83.085 35.655 83.255 35.825 ;
        RECT 83.545 35.655 83.715 35.825 ;
        RECT 84.005 35.655 84.175 35.825 ;
        RECT 84.465 35.655 84.635 35.825 ;
        RECT 84.925 35.655 85.095 35.825 ;
        RECT 85.385 35.655 85.555 35.825 ;
        RECT 85.845 35.655 86.015 35.825 ;
        RECT 86.305 35.655 86.475 35.825 ;
        RECT 86.765 35.655 86.935 35.825 ;
        RECT 87.225 35.655 87.395 35.825 ;
        RECT 87.685 35.655 87.855 35.825 ;
        RECT 88.145 35.655 88.315 35.825 ;
        RECT 88.605 35.655 88.775 35.825 ;
        RECT 89.065 35.655 89.235 35.825 ;
        RECT 89.525 35.655 89.695 35.825 ;
        RECT 89.985 35.655 90.155 35.825 ;
        RECT 90.445 35.655 90.615 35.825 ;
        RECT 90.905 35.655 91.075 35.825 ;
        RECT 91.365 35.655 91.535 35.825 ;
        RECT 91.825 35.655 91.995 35.825 ;
        RECT 92.285 35.655 92.455 35.825 ;
        RECT 92.745 35.655 92.915 35.825 ;
        RECT 93.205 35.655 93.375 35.825 ;
        RECT 93.665 35.655 93.835 35.825 ;
        RECT 94.125 35.655 94.295 35.825 ;
        RECT 94.585 35.655 94.755 35.825 ;
        RECT 95.045 35.655 95.215 35.825 ;
        RECT 95.505 35.655 95.675 35.825 ;
        RECT 95.965 35.655 96.135 35.825 ;
        RECT 96.425 35.655 96.595 35.825 ;
        RECT 96.885 35.655 97.055 35.825 ;
        RECT 97.345 35.655 97.515 35.825 ;
        RECT 97.805 35.655 97.975 35.825 ;
        RECT 98.265 35.655 98.435 35.825 ;
        RECT 98.725 35.655 98.895 35.825 ;
        RECT 99.185 35.655 99.355 35.825 ;
        RECT 99.645 35.655 99.815 35.825 ;
        RECT 16.845 30.215 17.015 30.385 ;
        RECT 17.305 30.215 17.475 30.385 ;
        RECT 17.765 30.215 17.935 30.385 ;
        RECT 18.225 30.215 18.395 30.385 ;
        RECT 18.685 30.215 18.855 30.385 ;
        RECT 19.145 30.215 19.315 30.385 ;
        RECT 19.605 30.215 19.775 30.385 ;
        RECT 20.065 30.215 20.235 30.385 ;
        RECT 20.525 30.215 20.695 30.385 ;
        RECT 20.985 30.215 21.155 30.385 ;
        RECT 21.445 30.215 21.615 30.385 ;
        RECT 21.905 30.215 22.075 30.385 ;
        RECT 22.365 30.215 22.535 30.385 ;
        RECT 22.825 30.215 22.995 30.385 ;
        RECT 23.285 30.215 23.455 30.385 ;
        RECT 23.745 30.215 23.915 30.385 ;
        RECT 24.205 30.215 24.375 30.385 ;
        RECT 24.665 30.215 24.835 30.385 ;
        RECT 25.125 30.215 25.295 30.385 ;
        RECT 25.585 30.215 25.755 30.385 ;
        RECT 26.045 30.215 26.215 30.385 ;
        RECT 26.505 30.215 26.675 30.385 ;
        RECT 26.965 30.215 27.135 30.385 ;
        RECT 27.425 30.215 27.595 30.385 ;
        RECT 27.885 30.215 28.055 30.385 ;
        RECT 28.345 30.215 28.515 30.385 ;
        RECT 28.805 30.215 28.975 30.385 ;
        RECT 29.265 30.215 29.435 30.385 ;
        RECT 29.725 30.215 29.895 30.385 ;
        RECT 30.185 30.215 30.355 30.385 ;
        RECT 30.645 30.215 30.815 30.385 ;
        RECT 31.105 30.215 31.275 30.385 ;
        RECT 31.565 30.215 31.735 30.385 ;
        RECT 32.025 30.215 32.195 30.385 ;
        RECT 32.485 30.215 32.655 30.385 ;
        RECT 32.945 30.215 33.115 30.385 ;
        RECT 33.405 30.215 33.575 30.385 ;
        RECT 33.865 30.215 34.035 30.385 ;
        RECT 34.325 30.215 34.495 30.385 ;
        RECT 34.785 30.215 34.955 30.385 ;
        RECT 35.245 30.215 35.415 30.385 ;
        RECT 35.705 30.215 35.875 30.385 ;
        RECT 36.165 30.215 36.335 30.385 ;
        RECT 36.625 30.215 36.795 30.385 ;
        RECT 37.085 30.215 37.255 30.385 ;
        RECT 37.545 30.215 37.715 30.385 ;
        RECT 38.005 30.215 38.175 30.385 ;
        RECT 38.465 30.215 38.635 30.385 ;
        RECT 38.925 30.215 39.095 30.385 ;
        RECT 39.385 30.215 39.555 30.385 ;
        RECT 39.845 30.215 40.015 30.385 ;
        RECT 40.305 30.215 40.475 30.385 ;
        RECT 40.765 30.215 40.935 30.385 ;
        RECT 41.225 30.215 41.395 30.385 ;
        RECT 41.685 30.215 41.855 30.385 ;
        RECT 42.145 30.215 42.315 30.385 ;
        RECT 42.605 30.215 42.775 30.385 ;
        RECT 43.065 30.215 43.235 30.385 ;
        RECT 43.525 30.215 43.695 30.385 ;
        RECT 43.985 30.215 44.155 30.385 ;
        RECT 44.445 30.215 44.615 30.385 ;
        RECT 44.905 30.215 45.075 30.385 ;
        RECT 45.365 30.215 45.535 30.385 ;
        RECT 45.825 30.215 45.995 30.385 ;
        RECT 46.285 30.215 46.455 30.385 ;
        RECT 46.745 30.215 46.915 30.385 ;
        RECT 47.205 30.215 47.375 30.385 ;
        RECT 47.665 30.215 47.835 30.385 ;
        RECT 48.125 30.215 48.295 30.385 ;
        RECT 48.585 30.215 48.755 30.385 ;
        RECT 49.045 30.215 49.215 30.385 ;
        RECT 49.505 30.215 49.675 30.385 ;
        RECT 49.965 30.215 50.135 30.385 ;
        RECT 50.425 30.215 50.595 30.385 ;
        RECT 50.885 30.215 51.055 30.385 ;
        RECT 51.345 30.215 51.515 30.385 ;
        RECT 51.805 30.215 51.975 30.385 ;
        RECT 52.265 30.215 52.435 30.385 ;
        RECT 52.725 30.215 52.895 30.385 ;
        RECT 53.185 30.215 53.355 30.385 ;
        RECT 53.645 30.215 53.815 30.385 ;
        RECT 54.105 30.215 54.275 30.385 ;
        RECT 54.565 30.215 54.735 30.385 ;
        RECT 55.025 30.215 55.195 30.385 ;
        RECT 55.485 30.215 55.655 30.385 ;
        RECT 55.945 30.215 56.115 30.385 ;
        RECT 56.405 30.215 56.575 30.385 ;
        RECT 56.865 30.215 57.035 30.385 ;
        RECT 57.325 30.215 57.495 30.385 ;
        RECT 57.785 30.215 57.955 30.385 ;
        RECT 58.245 30.215 58.415 30.385 ;
        RECT 58.705 30.215 58.875 30.385 ;
        RECT 59.165 30.215 59.335 30.385 ;
        RECT 59.625 30.215 59.795 30.385 ;
        RECT 60.085 30.215 60.255 30.385 ;
        RECT 60.545 30.215 60.715 30.385 ;
        RECT 61.005 30.215 61.175 30.385 ;
        RECT 61.465 30.215 61.635 30.385 ;
        RECT 61.925 30.215 62.095 30.385 ;
        RECT 62.385 30.215 62.555 30.385 ;
        RECT 62.845 30.215 63.015 30.385 ;
        RECT 63.305 30.215 63.475 30.385 ;
        RECT 63.765 30.215 63.935 30.385 ;
        RECT 64.225 30.215 64.395 30.385 ;
        RECT 64.685 30.215 64.855 30.385 ;
        RECT 65.145 30.215 65.315 30.385 ;
        RECT 65.605 30.215 65.775 30.385 ;
        RECT 66.065 30.215 66.235 30.385 ;
        RECT 66.525 30.215 66.695 30.385 ;
        RECT 66.985 30.215 67.155 30.385 ;
        RECT 67.445 30.215 67.615 30.385 ;
        RECT 67.905 30.215 68.075 30.385 ;
        RECT 68.365 30.215 68.535 30.385 ;
        RECT 68.825 30.215 68.995 30.385 ;
        RECT 69.285 30.215 69.455 30.385 ;
        RECT 69.745 30.215 69.915 30.385 ;
        RECT 70.205 30.215 70.375 30.385 ;
        RECT 70.665 30.215 70.835 30.385 ;
        RECT 71.125 30.215 71.295 30.385 ;
        RECT 71.585 30.215 71.755 30.385 ;
        RECT 72.045 30.215 72.215 30.385 ;
        RECT 72.505 30.215 72.675 30.385 ;
        RECT 72.965 30.215 73.135 30.385 ;
        RECT 73.425 30.215 73.595 30.385 ;
        RECT 73.885 30.215 74.055 30.385 ;
        RECT 74.345 30.215 74.515 30.385 ;
        RECT 74.805 30.215 74.975 30.385 ;
        RECT 75.265 30.215 75.435 30.385 ;
        RECT 75.725 30.215 75.895 30.385 ;
        RECT 76.185 30.215 76.355 30.385 ;
        RECT 76.645 30.215 76.815 30.385 ;
        RECT 77.105 30.215 77.275 30.385 ;
        RECT 77.565 30.215 77.735 30.385 ;
        RECT 78.025 30.215 78.195 30.385 ;
        RECT 78.485 30.215 78.655 30.385 ;
        RECT 78.945 30.215 79.115 30.385 ;
        RECT 79.405 30.215 79.575 30.385 ;
        RECT 79.865 30.215 80.035 30.385 ;
        RECT 80.325 30.215 80.495 30.385 ;
        RECT 80.785 30.215 80.955 30.385 ;
        RECT 81.245 30.215 81.415 30.385 ;
        RECT 81.705 30.215 81.875 30.385 ;
        RECT 82.165 30.215 82.335 30.385 ;
        RECT 82.625 30.215 82.795 30.385 ;
        RECT 83.085 30.215 83.255 30.385 ;
        RECT 83.545 30.215 83.715 30.385 ;
        RECT 84.005 30.215 84.175 30.385 ;
        RECT 84.465 30.215 84.635 30.385 ;
        RECT 84.925 30.215 85.095 30.385 ;
        RECT 85.385 30.215 85.555 30.385 ;
        RECT 85.845 30.215 86.015 30.385 ;
        RECT 86.305 30.215 86.475 30.385 ;
        RECT 86.765 30.215 86.935 30.385 ;
        RECT 87.225 30.215 87.395 30.385 ;
        RECT 87.685 30.215 87.855 30.385 ;
        RECT 88.145 30.215 88.315 30.385 ;
        RECT 88.605 30.215 88.775 30.385 ;
        RECT 89.065 30.215 89.235 30.385 ;
        RECT 89.525 30.215 89.695 30.385 ;
        RECT 89.985 30.215 90.155 30.385 ;
        RECT 90.445 30.215 90.615 30.385 ;
        RECT 90.905 30.215 91.075 30.385 ;
        RECT 91.365 30.215 91.535 30.385 ;
        RECT 91.825 30.215 91.995 30.385 ;
        RECT 92.285 30.215 92.455 30.385 ;
        RECT 92.745 30.215 92.915 30.385 ;
        RECT 93.205 30.215 93.375 30.385 ;
        RECT 93.665 30.215 93.835 30.385 ;
        RECT 94.125 30.215 94.295 30.385 ;
        RECT 94.585 30.215 94.755 30.385 ;
        RECT 95.045 30.215 95.215 30.385 ;
        RECT 95.505 30.215 95.675 30.385 ;
        RECT 95.965 30.215 96.135 30.385 ;
        RECT 96.425 30.215 96.595 30.385 ;
        RECT 96.885 30.215 97.055 30.385 ;
        RECT 97.345 30.215 97.515 30.385 ;
        RECT 97.805 30.215 97.975 30.385 ;
        RECT 98.265 30.215 98.435 30.385 ;
        RECT 98.725 30.215 98.895 30.385 ;
        RECT 99.185 30.215 99.355 30.385 ;
        RECT 99.645 30.215 99.815 30.385 ;
        RECT 16.845 24.775 17.015 24.945 ;
        RECT 17.305 24.775 17.475 24.945 ;
        RECT 17.765 24.775 17.935 24.945 ;
        RECT 18.225 24.775 18.395 24.945 ;
        RECT 18.685 24.775 18.855 24.945 ;
        RECT 19.145 24.775 19.315 24.945 ;
        RECT 19.605 24.775 19.775 24.945 ;
        RECT 20.065 24.775 20.235 24.945 ;
        RECT 20.525 24.775 20.695 24.945 ;
        RECT 20.985 24.775 21.155 24.945 ;
        RECT 21.445 24.775 21.615 24.945 ;
        RECT 21.905 24.775 22.075 24.945 ;
        RECT 22.365 24.775 22.535 24.945 ;
        RECT 22.825 24.775 22.995 24.945 ;
        RECT 23.285 24.775 23.455 24.945 ;
        RECT 23.745 24.775 23.915 24.945 ;
        RECT 24.205 24.775 24.375 24.945 ;
        RECT 24.665 24.775 24.835 24.945 ;
        RECT 25.125 24.775 25.295 24.945 ;
        RECT 25.585 24.775 25.755 24.945 ;
        RECT 26.045 24.775 26.215 24.945 ;
        RECT 26.505 24.775 26.675 24.945 ;
        RECT 26.965 24.775 27.135 24.945 ;
        RECT 27.425 24.775 27.595 24.945 ;
        RECT 27.885 24.775 28.055 24.945 ;
        RECT 28.345 24.775 28.515 24.945 ;
        RECT 28.805 24.775 28.975 24.945 ;
        RECT 29.265 24.775 29.435 24.945 ;
        RECT 29.725 24.775 29.895 24.945 ;
        RECT 30.185 24.775 30.355 24.945 ;
        RECT 30.645 24.775 30.815 24.945 ;
        RECT 31.105 24.775 31.275 24.945 ;
        RECT 31.565 24.775 31.735 24.945 ;
        RECT 32.025 24.775 32.195 24.945 ;
        RECT 32.485 24.775 32.655 24.945 ;
        RECT 32.945 24.775 33.115 24.945 ;
        RECT 33.405 24.775 33.575 24.945 ;
        RECT 33.865 24.775 34.035 24.945 ;
        RECT 34.325 24.775 34.495 24.945 ;
        RECT 34.785 24.775 34.955 24.945 ;
        RECT 35.245 24.775 35.415 24.945 ;
        RECT 35.705 24.775 35.875 24.945 ;
        RECT 36.165 24.775 36.335 24.945 ;
        RECT 36.625 24.775 36.795 24.945 ;
        RECT 37.085 24.775 37.255 24.945 ;
        RECT 37.545 24.775 37.715 24.945 ;
        RECT 38.005 24.775 38.175 24.945 ;
        RECT 38.465 24.775 38.635 24.945 ;
        RECT 38.925 24.775 39.095 24.945 ;
        RECT 39.385 24.775 39.555 24.945 ;
        RECT 39.845 24.775 40.015 24.945 ;
        RECT 40.305 24.775 40.475 24.945 ;
        RECT 40.765 24.775 40.935 24.945 ;
        RECT 41.225 24.775 41.395 24.945 ;
        RECT 41.685 24.775 41.855 24.945 ;
        RECT 42.145 24.775 42.315 24.945 ;
        RECT 42.605 24.775 42.775 24.945 ;
        RECT 43.065 24.775 43.235 24.945 ;
        RECT 43.525 24.775 43.695 24.945 ;
        RECT 43.985 24.775 44.155 24.945 ;
        RECT 44.445 24.775 44.615 24.945 ;
        RECT 44.905 24.775 45.075 24.945 ;
        RECT 45.365 24.775 45.535 24.945 ;
        RECT 45.825 24.775 45.995 24.945 ;
        RECT 46.285 24.775 46.455 24.945 ;
        RECT 46.745 24.775 46.915 24.945 ;
        RECT 47.205 24.775 47.375 24.945 ;
        RECT 47.665 24.775 47.835 24.945 ;
        RECT 48.125 24.775 48.295 24.945 ;
        RECT 48.585 24.775 48.755 24.945 ;
        RECT 49.045 24.775 49.215 24.945 ;
        RECT 49.505 24.775 49.675 24.945 ;
        RECT 49.965 24.775 50.135 24.945 ;
        RECT 50.425 24.775 50.595 24.945 ;
        RECT 50.885 24.775 51.055 24.945 ;
        RECT 51.345 24.775 51.515 24.945 ;
        RECT 51.805 24.775 51.975 24.945 ;
        RECT 52.265 24.775 52.435 24.945 ;
        RECT 52.725 24.775 52.895 24.945 ;
        RECT 53.185 24.775 53.355 24.945 ;
        RECT 53.645 24.775 53.815 24.945 ;
        RECT 54.105 24.775 54.275 24.945 ;
        RECT 54.565 24.775 54.735 24.945 ;
        RECT 55.025 24.775 55.195 24.945 ;
        RECT 55.485 24.775 55.655 24.945 ;
        RECT 55.945 24.775 56.115 24.945 ;
        RECT 56.405 24.775 56.575 24.945 ;
        RECT 56.865 24.775 57.035 24.945 ;
        RECT 57.325 24.775 57.495 24.945 ;
        RECT 57.785 24.775 57.955 24.945 ;
        RECT 58.245 24.775 58.415 24.945 ;
        RECT 58.705 24.775 58.875 24.945 ;
        RECT 59.165 24.775 59.335 24.945 ;
        RECT 59.625 24.775 59.795 24.945 ;
        RECT 60.085 24.775 60.255 24.945 ;
        RECT 60.545 24.775 60.715 24.945 ;
        RECT 61.005 24.775 61.175 24.945 ;
        RECT 61.465 24.775 61.635 24.945 ;
        RECT 61.925 24.775 62.095 24.945 ;
        RECT 62.385 24.775 62.555 24.945 ;
        RECT 62.845 24.775 63.015 24.945 ;
        RECT 63.305 24.775 63.475 24.945 ;
        RECT 63.765 24.775 63.935 24.945 ;
        RECT 64.225 24.775 64.395 24.945 ;
        RECT 64.685 24.775 64.855 24.945 ;
        RECT 65.145 24.775 65.315 24.945 ;
        RECT 65.605 24.775 65.775 24.945 ;
        RECT 66.065 24.775 66.235 24.945 ;
        RECT 66.525 24.775 66.695 24.945 ;
        RECT 66.985 24.775 67.155 24.945 ;
        RECT 67.445 24.775 67.615 24.945 ;
        RECT 67.905 24.775 68.075 24.945 ;
        RECT 68.365 24.775 68.535 24.945 ;
        RECT 68.825 24.775 68.995 24.945 ;
        RECT 69.285 24.775 69.455 24.945 ;
        RECT 69.745 24.775 69.915 24.945 ;
        RECT 70.205 24.775 70.375 24.945 ;
        RECT 70.665 24.775 70.835 24.945 ;
        RECT 71.125 24.775 71.295 24.945 ;
        RECT 71.585 24.775 71.755 24.945 ;
        RECT 72.045 24.775 72.215 24.945 ;
        RECT 72.505 24.775 72.675 24.945 ;
        RECT 72.965 24.775 73.135 24.945 ;
        RECT 73.425 24.775 73.595 24.945 ;
        RECT 73.885 24.775 74.055 24.945 ;
        RECT 74.345 24.775 74.515 24.945 ;
        RECT 74.805 24.775 74.975 24.945 ;
        RECT 75.265 24.775 75.435 24.945 ;
        RECT 75.725 24.775 75.895 24.945 ;
        RECT 76.185 24.775 76.355 24.945 ;
        RECT 76.645 24.775 76.815 24.945 ;
        RECT 77.105 24.775 77.275 24.945 ;
        RECT 77.565 24.775 77.735 24.945 ;
        RECT 78.025 24.775 78.195 24.945 ;
        RECT 78.485 24.775 78.655 24.945 ;
        RECT 78.945 24.775 79.115 24.945 ;
        RECT 79.405 24.775 79.575 24.945 ;
        RECT 79.865 24.775 80.035 24.945 ;
        RECT 80.325 24.775 80.495 24.945 ;
        RECT 80.785 24.775 80.955 24.945 ;
        RECT 81.245 24.775 81.415 24.945 ;
        RECT 81.705 24.775 81.875 24.945 ;
        RECT 82.165 24.775 82.335 24.945 ;
        RECT 82.625 24.775 82.795 24.945 ;
        RECT 83.085 24.775 83.255 24.945 ;
        RECT 83.545 24.775 83.715 24.945 ;
        RECT 84.005 24.775 84.175 24.945 ;
        RECT 84.465 24.775 84.635 24.945 ;
        RECT 84.925 24.775 85.095 24.945 ;
        RECT 85.385 24.775 85.555 24.945 ;
        RECT 85.845 24.775 86.015 24.945 ;
        RECT 86.305 24.775 86.475 24.945 ;
        RECT 86.765 24.775 86.935 24.945 ;
        RECT 87.225 24.775 87.395 24.945 ;
        RECT 87.685 24.775 87.855 24.945 ;
        RECT 88.145 24.775 88.315 24.945 ;
        RECT 88.605 24.775 88.775 24.945 ;
        RECT 89.065 24.775 89.235 24.945 ;
        RECT 89.525 24.775 89.695 24.945 ;
        RECT 89.985 24.775 90.155 24.945 ;
        RECT 90.445 24.775 90.615 24.945 ;
        RECT 90.905 24.775 91.075 24.945 ;
        RECT 91.365 24.775 91.535 24.945 ;
        RECT 91.825 24.775 91.995 24.945 ;
        RECT 92.285 24.775 92.455 24.945 ;
        RECT 92.745 24.775 92.915 24.945 ;
        RECT 93.205 24.775 93.375 24.945 ;
        RECT 93.665 24.775 93.835 24.945 ;
        RECT 94.125 24.775 94.295 24.945 ;
        RECT 94.585 24.775 94.755 24.945 ;
        RECT 95.045 24.775 95.215 24.945 ;
        RECT 95.505 24.775 95.675 24.945 ;
        RECT 95.965 24.775 96.135 24.945 ;
        RECT 96.425 24.775 96.595 24.945 ;
        RECT 96.885 24.775 97.055 24.945 ;
        RECT 97.345 24.775 97.515 24.945 ;
        RECT 97.805 24.775 97.975 24.945 ;
        RECT 98.265 24.775 98.435 24.945 ;
        RECT 98.725 24.775 98.895 24.945 ;
        RECT 99.185 24.775 99.355 24.945 ;
        RECT 99.645 24.775 99.815 24.945 ;
        RECT 16.845 19.335 17.015 19.505 ;
        RECT 17.305 19.335 17.475 19.505 ;
        RECT 17.765 19.335 17.935 19.505 ;
        RECT 18.225 19.335 18.395 19.505 ;
        RECT 18.685 19.335 18.855 19.505 ;
        RECT 19.145 19.335 19.315 19.505 ;
        RECT 19.605 19.335 19.775 19.505 ;
        RECT 20.065 19.335 20.235 19.505 ;
        RECT 20.525 19.335 20.695 19.505 ;
        RECT 20.985 19.335 21.155 19.505 ;
        RECT 21.445 19.335 21.615 19.505 ;
        RECT 21.905 19.335 22.075 19.505 ;
        RECT 22.365 19.335 22.535 19.505 ;
        RECT 22.825 19.335 22.995 19.505 ;
        RECT 23.285 19.335 23.455 19.505 ;
        RECT 23.745 19.335 23.915 19.505 ;
        RECT 24.205 19.335 24.375 19.505 ;
        RECT 24.665 19.335 24.835 19.505 ;
        RECT 25.125 19.335 25.295 19.505 ;
        RECT 25.585 19.335 25.755 19.505 ;
        RECT 26.045 19.335 26.215 19.505 ;
        RECT 26.505 19.335 26.675 19.505 ;
        RECT 26.965 19.335 27.135 19.505 ;
        RECT 27.425 19.335 27.595 19.505 ;
        RECT 27.885 19.335 28.055 19.505 ;
        RECT 28.345 19.335 28.515 19.505 ;
        RECT 28.805 19.335 28.975 19.505 ;
        RECT 29.265 19.335 29.435 19.505 ;
        RECT 29.725 19.335 29.895 19.505 ;
        RECT 30.185 19.335 30.355 19.505 ;
        RECT 30.645 19.335 30.815 19.505 ;
        RECT 31.105 19.335 31.275 19.505 ;
        RECT 31.565 19.335 31.735 19.505 ;
        RECT 32.025 19.335 32.195 19.505 ;
        RECT 32.485 19.335 32.655 19.505 ;
        RECT 32.945 19.335 33.115 19.505 ;
        RECT 33.405 19.335 33.575 19.505 ;
        RECT 33.865 19.335 34.035 19.505 ;
        RECT 34.325 19.335 34.495 19.505 ;
        RECT 34.785 19.335 34.955 19.505 ;
        RECT 35.245 19.335 35.415 19.505 ;
        RECT 35.705 19.335 35.875 19.505 ;
        RECT 36.165 19.335 36.335 19.505 ;
        RECT 36.625 19.335 36.795 19.505 ;
        RECT 37.085 19.335 37.255 19.505 ;
        RECT 37.545 19.335 37.715 19.505 ;
        RECT 38.005 19.335 38.175 19.505 ;
        RECT 38.465 19.335 38.635 19.505 ;
        RECT 38.925 19.335 39.095 19.505 ;
        RECT 39.385 19.335 39.555 19.505 ;
        RECT 39.845 19.335 40.015 19.505 ;
        RECT 40.305 19.335 40.475 19.505 ;
        RECT 40.765 19.335 40.935 19.505 ;
        RECT 41.225 19.335 41.395 19.505 ;
        RECT 41.685 19.335 41.855 19.505 ;
        RECT 42.145 19.335 42.315 19.505 ;
        RECT 42.605 19.335 42.775 19.505 ;
        RECT 43.065 19.335 43.235 19.505 ;
        RECT 43.525 19.335 43.695 19.505 ;
        RECT 43.985 19.335 44.155 19.505 ;
        RECT 44.445 19.335 44.615 19.505 ;
        RECT 44.905 19.335 45.075 19.505 ;
        RECT 45.365 19.335 45.535 19.505 ;
        RECT 45.825 19.335 45.995 19.505 ;
        RECT 46.285 19.335 46.455 19.505 ;
        RECT 46.745 19.335 46.915 19.505 ;
        RECT 47.205 19.335 47.375 19.505 ;
        RECT 47.665 19.335 47.835 19.505 ;
        RECT 48.125 19.335 48.295 19.505 ;
        RECT 48.585 19.335 48.755 19.505 ;
        RECT 49.045 19.335 49.215 19.505 ;
        RECT 49.505 19.335 49.675 19.505 ;
        RECT 49.965 19.335 50.135 19.505 ;
        RECT 50.425 19.335 50.595 19.505 ;
        RECT 50.885 19.335 51.055 19.505 ;
        RECT 51.345 19.335 51.515 19.505 ;
        RECT 51.805 19.335 51.975 19.505 ;
        RECT 52.265 19.335 52.435 19.505 ;
        RECT 52.725 19.335 52.895 19.505 ;
        RECT 53.185 19.335 53.355 19.505 ;
        RECT 53.645 19.335 53.815 19.505 ;
        RECT 54.105 19.335 54.275 19.505 ;
        RECT 54.565 19.335 54.735 19.505 ;
        RECT 55.025 19.335 55.195 19.505 ;
        RECT 55.485 19.335 55.655 19.505 ;
        RECT 55.945 19.335 56.115 19.505 ;
        RECT 56.405 19.335 56.575 19.505 ;
        RECT 56.865 19.335 57.035 19.505 ;
        RECT 57.325 19.335 57.495 19.505 ;
        RECT 57.785 19.335 57.955 19.505 ;
        RECT 58.245 19.335 58.415 19.505 ;
        RECT 58.705 19.335 58.875 19.505 ;
        RECT 59.165 19.335 59.335 19.505 ;
        RECT 59.625 19.335 59.795 19.505 ;
        RECT 60.085 19.335 60.255 19.505 ;
        RECT 60.545 19.335 60.715 19.505 ;
        RECT 61.005 19.335 61.175 19.505 ;
        RECT 61.465 19.335 61.635 19.505 ;
        RECT 61.925 19.335 62.095 19.505 ;
        RECT 62.385 19.335 62.555 19.505 ;
        RECT 62.845 19.335 63.015 19.505 ;
        RECT 63.305 19.335 63.475 19.505 ;
        RECT 63.765 19.335 63.935 19.505 ;
        RECT 64.225 19.335 64.395 19.505 ;
        RECT 64.685 19.335 64.855 19.505 ;
        RECT 65.145 19.335 65.315 19.505 ;
        RECT 65.605 19.335 65.775 19.505 ;
        RECT 66.065 19.335 66.235 19.505 ;
        RECT 66.525 19.335 66.695 19.505 ;
        RECT 66.985 19.335 67.155 19.505 ;
        RECT 67.445 19.335 67.615 19.505 ;
        RECT 67.905 19.335 68.075 19.505 ;
        RECT 68.365 19.335 68.535 19.505 ;
        RECT 68.825 19.335 68.995 19.505 ;
        RECT 69.285 19.335 69.455 19.505 ;
        RECT 69.745 19.335 69.915 19.505 ;
        RECT 70.205 19.335 70.375 19.505 ;
        RECT 70.665 19.335 70.835 19.505 ;
        RECT 71.125 19.335 71.295 19.505 ;
        RECT 71.585 19.335 71.755 19.505 ;
        RECT 72.045 19.335 72.215 19.505 ;
        RECT 72.505 19.335 72.675 19.505 ;
        RECT 72.965 19.335 73.135 19.505 ;
        RECT 73.425 19.335 73.595 19.505 ;
        RECT 73.885 19.335 74.055 19.505 ;
        RECT 74.345 19.335 74.515 19.505 ;
        RECT 74.805 19.335 74.975 19.505 ;
        RECT 75.265 19.335 75.435 19.505 ;
        RECT 75.725 19.335 75.895 19.505 ;
        RECT 76.185 19.335 76.355 19.505 ;
        RECT 76.645 19.335 76.815 19.505 ;
        RECT 77.105 19.335 77.275 19.505 ;
        RECT 77.565 19.335 77.735 19.505 ;
        RECT 78.025 19.335 78.195 19.505 ;
        RECT 78.485 19.335 78.655 19.505 ;
        RECT 78.945 19.335 79.115 19.505 ;
        RECT 79.405 19.335 79.575 19.505 ;
        RECT 79.865 19.335 80.035 19.505 ;
        RECT 80.325 19.335 80.495 19.505 ;
        RECT 80.785 19.335 80.955 19.505 ;
        RECT 81.245 19.335 81.415 19.505 ;
        RECT 81.705 19.335 81.875 19.505 ;
        RECT 82.165 19.335 82.335 19.505 ;
        RECT 82.625 19.335 82.795 19.505 ;
        RECT 83.085 19.335 83.255 19.505 ;
        RECT 83.545 19.335 83.715 19.505 ;
        RECT 84.005 19.335 84.175 19.505 ;
        RECT 84.465 19.335 84.635 19.505 ;
        RECT 84.925 19.335 85.095 19.505 ;
        RECT 85.385 19.335 85.555 19.505 ;
        RECT 85.845 19.335 86.015 19.505 ;
        RECT 86.305 19.335 86.475 19.505 ;
        RECT 86.765 19.335 86.935 19.505 ;
        RECT 87.225 19.335 87.395 19.505 ;
        RECT 87.685 19.335 87.855 19.505 ;
        RECT 88.145 19.335 88.315 19.505 ;
        RECT 88.605 19.335 88.775 19.505 ;
        RECT 89.065 19.335 89.235 19.505 ;
        RECT 89.525 19.335 89.695 19.505 ;
        RECT 89.985 19.335 90.155 19.505 ;
        RECT 90.445 19.335 90.615 19.505 ;
        RECT 90.905 19.335 91.075 19.505 ;
        RECT 91.365 19.335 91.535 19.505 ;
        RECT 91.825 19.335 91.995 19.505 ;
        RECT 92.285 19.335 92.455 19.505 ;
        RECT 92.745 19.335 92.915 19.505 ;
        RECT 93.205 19.335 93.375 19.505 ;
        RECT 93.665 19.335 93.835 19.505 ;
        RECT 94.125 19.335 94.295 19.505 ;
        RECT 94.585 19.335 94.755 19.505 ;
        RECT 95.045 19.335 95.215 19.505 ;
        RECT 95.505 19.335 95.675 19.505 ;
        RECT 95.965 19.335 96.135 19.505 ;
        RECT 96.425 19.335 96.595 19.505 ;
        RECT 96.885 19.335 97.055 19.505 ;
        RECT 97.345 19.335 97.515 19.505 ;
        RECT 97.805 19.335 97.975 19.505 ;
        RECT 98.265 19.335 98.435 19.505 ;
        RECT 98.725 19.335 98.895 19.505 ;
        RECT 99.185 19.335 99.355 19.505 ;
        RECT 99.645 19.335 99.815 19.505 ;
      LAYER met1 ;
        RECT 16.700 95.340 99.960 95.820 ;
        RECT 16.700 89.900 99.960 90.380 ;
        RECT 16.700 84.460 99.960 84.940 ;
        RECT 16.700 79.020 99.960 79.500 ;
        RECT 16.700 73.580 99.960 74.060 ;
        RECT 16.700 68.140 99.960 68.620 ;
        RECT 16.700 62.700 99.960 63.180 ;
        RECT 16.700 57.260 99.960 57.740 ;
        RECT 16.700 51.820 99.960 52.300 ;
        RECT 16.700 46.380 99.960 46.860 ;
        RECT 16.700 40.940 99.960 41.420 ;
        RECT 16.700 35.500 99.960 35.980 ;
        RECT 16.700 30.060 99.960 30.540 ;
        RECT 16.700 24.620 99.960 25.100 ;
        RECT 16.700 19.180 99.960 19.660 ;
      LAYER via ;
        RECT 43.840 95.450 44.100 95.710 ;
        RECT 44.160 95.450 44.420 95.710 ;
        RECT 44.480 95.450 44.740 95.710 ;
        RECT 44.800 95.450 45.060 95.710 ;
        RECT 71.595 95.450 71.855 95.710 ;
        RECT 71.915 95.450 72.175 95.710 ;
        RECT 72.235 95.450 72.495 95.710 ;
        RECT 72.555 95.450 72.815 95.710 ;
        RECT 43.840 90.010 44.100 90.270 ;
        RECT 44.160 90.010 44.420 90.270 ;
        RECT 44.480 90.010 44.740 90.270 ;
        RECT 44.800 90.010 45.060 90.270 ;
        RECT 71.595 90.010 71.855 90.270 ;
        RECT 71.915 90.010 72.175 90.270 ;
        RECT 72.235 90.010 72.495 90.270 ;
        RECT 72.555 90.010 72.815 90.270 ;
        RECT 43.840 84.570 44.100 84.830 ;
        RECT 44.160 84.570 44.420 84.830 ;
        RECT 44.480 84.570 44.740 84.830 ;
        RECT 44.800 84.570 45.060 84.830 ;
        RECT 71.595 84.570 71.855 84.830 ;
        RECT 71.915 84.570 72.175 84.830 ;
        RECT 72.235 84.570 72.495 84.830 ;
        RECT 72.555 84.570 72.815 84.830 ;
        RECT 43.840 79.130 44.100 79.390 ;
        RECT 44.160 79.130 44.420 79.390 ;
        RECT 44.480 79.130 44.740 79.390 ;
        RECT 44.800 79.130 45.060 79.390 ;
        RECT 71.595 79.130 71.855 79.390 ;
        RECT 71.915 79.130 72.175 79.390 ;
        RECT 72.235 79.130 72.495 79.390 ;
        RECT 72.555 79.130 72.815 79.390 ;
        RECT 43.840 73.690 44.100 73.950 ;
        RECT 44.160 73.690 44.420 73.950 ;
        RECT 44.480 73.690 44.740 73.950 ;
        RECT 44.800 73.690 45.060 73.950 ;
        RECT 71.595 73.690 71.855 73.950 ;
        RECT 71.915 73.690 72.175 73.950 ;
        RECT 72.235 73.690 72.495 73.950 ;
        RECT 72.555 73.690 72.815 73.950 ;
        RECT 43.840 68.250 44.100 68.510 ;
        RECT 44.160 68.250 44.420 68.510 ;
        RECT 44.480 68.250 44.740 68.510 ;
        RECT 44.800 68.250 45.060 68.510 ;
        RECT 71.595 68.250 71.855 68.510 ;
        RECT 71.915 68.250 72.175 68.510 ;
        RECT 72.235 68.250 72.495 68.510 ;
        RECT 72.555 68.250 72.815 68.510 ;
        RECT 43.840 62.810 44.100 63.070 ;
        RECT 44.160 62.810 44.420 63.070 ;
        RECT 44.480 62.810 44.740 63.070 ;
        RECT 44.800 62.810 45.060 63.070 ;
        RECT 71.595 62.810 71.855 63.070 ;
        RECT 71.915 62.810 72.175 63.070 ;
        RECT 72.235 62.810 72.495 63.070 ;
        RECT 72.555 62.810 72.815 63.070 ;
        RECT 43.840 57.370 44.100 57.630 ;
        RECT 44.160 57.370 44.420 57.630 ;
        RECT 44.480 57.370 44.740 57.630 ;
        RECT 44.800 57.370 45.060 57.630 ;
        RECT 71.595 57.370 71.855 57.630 ;
        RECT 71.915 57.370 72.175 57.630 ;
        RECT 72.235 57.370 72.495 57.630 ;
        RECT 72.555 57.370 72.815 57.630 ;
        RECT 43.840 51.930 44.100 52.190 ;
        RECT 44.160 51.930 44.420 52.190 ;
        RECT 44.480 51.930 44.740 52.190 ;
        RECT 44.800 51.930 45.060 52.190 ;
        RECT 71.595 51.930 71.855 52.190 ;
        RECT 71.915 51.930 72.175 52.190 ;
        RECT 72.235 51.930 72.495 52.190 ;
        RECT 72.555 51.930 72.815 52.190 ;
        RECT 43.840 46.490 44.100 46.750 ;
        RECT 44.160 46.490 44.420 46.750 ;
        RECT 44.480 46.490 44.740 46.750 ;
        RECT 44.800 46.490 45.060 46.750 ;
        RECT 71.595 46.490 71.855 46.750 ;
        RECT 71.915 46.490 72.175 46.750 ;
        RECT 72.235 46.490 72.495 46.750 ;
        RECT 72.555 46.490 72.815 46.750 ;
        RECT 43.840 41.050 44.100 41.310 ;
        RECT 44.160 41.050 44.420 41.310 ;
        RECT 44.480 41.050 44.740 41.310 ;
        RECT 44.800 41.050 45.060 41.310 ;
        RECT 71.595 41.050 71.855 41.310 ;
        RECT 71.915 41.050 72.175 41.310 ;
        RECT 72.235 41.050 72.495 41.310 ;
        RECT 72.555 41.050 72.815 41.310 ;
        RECT 43.840 35.610 44.100 35.870 ;
        RECT 44.160 35.610 44.420 35.870 ;
        RECT 44.480 35.610 44.740 35.870 ;
        RECT 44.800 35.610 45.060 35.870 ;
        RECT 71.595 35.610 71.855 35.870 ;
        RECT 71.915 35.610 72.175 35.870 ;
        RECT 72.235 35.610 72.495 35.870 ;
        RECT 72.555 35.610 72.815 35.870 ;
        RECT 43.840 30.170 44.100 30.430 ;
        RECT 44.160 30.170 44.420 30.430 ;
        RECT 44.480 30.170 44.740 30.430 ;
        RECT 44.800 30.170 45.060 30.430 ;
        RECT 71.595 30.170 71.855 30.430 ;
        RECT 71.915 30.170 72.175 30.430 ;
        RECT 72.235 30.170 72.495 30.430 ;
        RECT 72.555 30.170 72.815 30.430 ;
        RECT 43.840 24.730 44.100 24.990 ;
        RECT 44.160 24.730 44.420 24.990 ;
        RECT 44.480 24.730 44.740 24.990 ;
        RECT 44.800 24.730 45.060 24.990 ;
        RECT 71.595 24.730 71.855 24.990 ;
        RECT 71.915 24.730 72.175 24.990 ;
        RECT 72.235 24.730 72.495 24.990 ;
        RECT 72.555 24.730 72.815 24.990 ;
        RECT 43.840 19.290 44.100 19.550 ;
        RECT 44.160 19.290 44.420 19.550 ;
        RECT 44.480 19.290 44.740 19.550 ;
        RECT 44.800 19.290 45.060 19.550 ;
        RECT 71.595 19.290 71.855 19.550 ;
        RECT 71.915 19.290 72.175 19.550 ;
        RECT 72.235 19.290 72.495 19.550 ;
        RECT 72.555 19.290 72.815 19.550 ;
      LAYER met2 ;
        RECT 43.710 95.340 45.190 95.820 ;
        RECT 71.465 95.340 72.945 95.820 ;
        RECT 43.710 89.900 45.190 90.380 ;
        RECT 71.465 89.900 72.945 90.380 ;
        RECT 43.710 84.460 45.190 84.940 ;
        RECT 71.465 84.460 72.945 84.940 ;
        RECT 43.710 79.020 45.190 79.500 ;
        RECT 71.465 79.020 72.945 79.500 ;
        RECT 43.710 73.580 45.190 74.060 ;
        RECT 71.465 73.580 72.945 74.060 ;
        RECT 43.710 68.140 45.190 68.620 ;
        RECT 71.465 68.140 72.945 68.620 ;
        RECT 43.710 62.700 45.190 63.180 ;
        RECT 71.465 62.700 72.945 63.180 ;
        RECT 43.710 57.260 45.190 57.740 ;
        RECT 71.465 57.260 72.945 57.740 ;
        RECT 43.710 51.820 45.190 52.300 ;
        RECT 71.465 51.820 72.945 52.300 ;
        RECT 43.710 46.380 45.190 46.860 ;
        RECT 71.465 46.380 72.945 46.860 ;
        RECT 43.710 40.940 45.190 41.420 ;
        RECT 71.465 40.940 72.945 41.420 ;
        RECT 43.710 35.500 45.190 35.980 ;
        RECT 71.465 35.500 72.945 35.980 ;
        RECT 43.710 30.060 45.190 30.540 ;
        RECT 71.465 30.060 72.945 30.540 ;
        RECT 43.710 24.620 45.190 25.100 ;
        RECT 71.465 24.620 72.945 25.100 ;
        RECT 43.710 19.180 45.190 19.660 ;
        RECT 71.465 19.180 72.945 19.660 ;
      LAYER via2 ;
        RECT 43.710 95.440 43.990 95.720 ;
        RECT 44.110 95.440 44.390 95.720 ;
        RECT 44.510 95.440 44.790 95.720 ;
        RECT 44.910 95.440 45.190 95.720 ;
        RECT 71.465 95.440 71.745 95.720 ;
        RECT 71.865 95.440 72.145 95.720 ;
        RECT 72.265 95.440 72.545 95.720 ;
        RECT 72.665 95.440 72.945 95.720 ;
        RECT 43.710 90.000 43.990 90.280 ;
        RECT 44.110 90.000 44.390 90.280 ;
        RECT 44.510 90.000 44.790 90.280 ;
        RECT 44.910 90.000 45.190 90.280 ;
        RECT 71.465 90.000 71.745 90.280 ;
        RECT 71.865 90.000 72.145 90.280 ;
        RECT 72.265 90.000 72.545 90.280 ;
        RECT 72.665 90.000 72.945 90.280 ;
        RECT 43.710 84.560 43.990 84.840 ;
        RECT 44.110 84.560 44.390 84.840 ;
        RECT 44.510 84.560 44.790 84.840 ;
        RECT 44.910 84.560 45.190 84.840 ;
        RECT 71.465 84.560 71.745 84.840 ;
        RECT 71.865 84.560 72.145 84.840 ;
        RECT 72.265 84.560 72.545 84.840 ;
        RECT 72.665 84.560 72.945 84.840 ;
        RECT 43.710 79.120 43.990 79.400 ;
        RECT 44.110 79.120 44.390 79.400 ;
        RECT 44.510 79.120 44.790 79.400 ;
        RECT 44.910 79.120 45.190 79.400 ;
        RECT 71.465 79.120 71.745 79.400 ;
        RECT 71.865 79.120 72.145 79.400 ;
        RECT 72.265 79.120 72.545 79.400 ;
        RECT 72.665 79.120 72.945 79.400 ;
        RECT 43.710 73.680 43.990 73.960 ;
        RECT 44.110 73.680 44.390 73.960 ;
        RECT 44.510 73.680 44.790 73.960 ;
        RECT 44.910 73.680 45.190 73.960 ;
        RECT 71.465 73.680 71.745 73.960 ;
        RECT 71.865 73.680 72.145 73.960 ;
        RECT 72.265 73.680 72.545 73.960 ;
        RECT 72.665 73.680 72.945 73.960 ;
        RECT 43.710 68.240 43.990 68.520 ;
        RECT 44.110 68.240 44.390 68.520 ;
        RECT 44.510 68.240 44.790 68.520 ;
        RECT 44.910 68.240 45.190 68.520 ;
        RECT 71.465 68.240 71.745 68.520 ;
        RECT 71.865 68.240 72.145 68.520 ;
        RECT 72.265 68.240 72.545 68.520 ;
        RECT 72.665 68.240 72.945 68.520 ;
        RECT 43.710 62.800 43.990 63.080 ;
        RECT 44.110 62.800 44.390 63.080 ;
        RECT 44.510 62.800 44.790 63.080 ;
        RECT 44.910 62.800 45.190 63.080 ;
        RECT 71.465 62.800 71.745 63.080 ;
        RECT 71.865 62.800 72.145 63.080 ;
        RECT 72.265 62.800 72.545 63.080 ;
        RECT 72.665 62.800 72.945 63.080 ;
        RECT 43.710 57.360 43.990 57.640 ;
        RECT 44.110 57.360 44.390 57.640 ;
        RECT 44.510 57.360 44.790 57.640 ;
        RECT 44.910 57.360 45.190 57.640 ;
        RECT 71.465 57.360 71.745 57.640 ;
        RECT 71.865 57.360 72.145 57.640 ;
        RECT 72.265 57.360 72.545 57.640 ;
        RECT 72.665 57.360 72.945 57.640 ;
        RECT 43.710 51.920 43.990 52.200 ;
        RECT 44.110 51.920 44.390 52.200 ;
        RECT 44.510 51.920 44.790 52.200 ;
        RECT 44.910 51.920 45.190 52.200 ;
        RECT 71.465 51.920 71.745 52.200 ;
        RECT 71.865 51.920 72.145 52.200 ;
        RECT 72.265 51.920 72.545 52.200 ;
        RECT 72.665 51.920 72.945 52.200 ;
        RECT 43.710 46.480 43.990 46.760 ;
        RECT 44.110 46.480 44.390 46.760 ;
        RECT 44.510 46.480 44.790 46.760 ;
        RECT 44.910 46.480 45.190 46.760 ;
        RECT 71.465 46.480 71.745 46.760 ;
        RECT 71.865 46.480 72.145 46.760 ;
        RECT 72.265 46.480 72.545 46.760 ;
        RECT 72.665 46.480 72.945 46.760 ;
        RECT 43.710 41.040 43.990 41.320 ;
        RECT 44.110 41.040 44.390 41.320 ;
        RECT 44.510 41.040 44.790 41.320 ;
        RECT 44.910 41.040 45.190 41.320 ;
        RECT 71.465 41.040 71.745 41.320 ;
        RECT 71.865 41.040 72.145 41.320 ;
        RECT 72.265 41.040 72.545 41.320 ;
        RECT 72.665 41.040 72.945 41.320 ;
        RECT 43.710 35.600 43.990 35.880 ;
        RECT 44.110 35.600 44.390 35.880 ;
        RECT 44.510 35.600 44.790 35.880 ;
        RECT 44.910 35.600 45.190 35.880 ;
        RECT 71.465 35.600 71.745 35.880 ;
        RECT 71.865 35.600 72.145 35.880 ;
        RECT 72.265 35.600 72.545 35.880 ;
        RECT 72.665 35.600 72.945 35.880 ;
        RECT 43.710 30.160 43.990 30.440 ;
        RECT 44.110 30.160 44.390 30.440 ;
        RECT 44.510 30.160 44.790 30.440 ;
        RECT 44.910 30.160 45.190 30.440 ;
        RECT 71.465 30.160 71.745 30.440 ;
        RECT 71.865 30.160 72.145 30.440 ;
        RECT 72.265 30.160 72.545 30.440 ;
        RECT 72.665 30.160 72.945 30.440 ;
        RECT 43.710 24.720 43.990 25.000 ;
        RECT 44.110 24.720 44.390 25.000 ;
        RECT 44.510 24.720 44.790 25.000 ;
        RECT 44.910 24.720 45.190 25.000 ;
        RECT 71.465 24.720 71.745 25.000 ;
        RECT 71.865 24.720 72.145 25.000 ;
        RECT 72.265 24.720 72.545 25.000 ;
        RECT 72.665 24.720 72.945 25.000 ;
        RECT 43.710 19.280 43.990 19.560 ;
        RECT 44.110 19.280 44.390 19.560 ;
        RECT 44.510 19.280 44.790 19.560 ;
        RECT 44.910 19.280 45.190 19.560 ;
        RECT 71.465 19.280 71.745 19.560 ;
        RECT 71.865 19.280 72.145 19.560 ;
        RECT 72.265 19.280 72.545 19.560 ;
        RECT 72.665 19.280 72.945 19.560 ;
      LAYER met3 ;
        RECT 43.650 95.415 45.250 95.745 ;
        RECT 71.405 95.415 73.005 95.745 ;
        RECT 43.650 89.975 45.250 90.305 ;
        RECT 71.405 89.975 73.005 90.305 ;
        RECT 43.650 84.535 45.250 84.865 ;
        RECT 71.405 84.535 73.005 84.865 ;
        RECT 43.650 79.095 45.250 79.425 ;
        RECT 71.405 79.095 73.005 79.425 ;
        RECT 43.650 73.655 45.250 73.985 ;
        RECT 71.405 73.655 73.005 73.985 ;
        RECT 43.650 68.215 45.250 68.545 ;
        RECT 71.405 68.215 73.005 68.545 ;
        RECT 43.650 62.775 45.250 63.105 ;
        RECT 71.405 62.775 73.005 63.105 ;
        RECT 43.650 57.335 45.250 57.665 ;
        RECT 71.405 57.335 73.005 57.665 ;
        RECT 43.650 51.895 45.250 52.225 ;
        RECT 71.405 51.895 73.005 52.225 ;
        RECT 43.650 46.455 45.250 46.785 ;
        RECT 71.405 46.455 73.005 46.785 ;
        RECT 43.650 41.015 45.250 41.345 ;
        RECT 71.405 41.015 73.005 41.345 ;
        RECT 43.650 35.575 45.250 35.905 ;
        RECT 71.405 35.575 73.005 35.905 ;
        RECT 43.650 30.135 45.250 30.465 ;
        RECT 71.405 30.135 73.005 30.465 ;
        RECT 43.650 24.695 45.250 25.025 ;
        RECT 71.405 24.695 73.005 25.025 ;
        RECT 43.650 19.255 45.250 19.585 ;
        RECT 71.405 19.255 73.005 19.585 ;
      LAYER via3 ;
        RECT 43.690 95.420 44.010 95.740 ;
        RECT 44.090 95.420 44.410 95.740 ;
        RECT 44.490 95.420 44.810 95.740 ;
        RECT 44.890 95.420 45.210 95.740 ;
        RECT 71.445 95.420 71.765 95.740 ;
        RECT 71.845 95.420 72.165 95.740 ;
        RECT 72.245 95.420 72.565 95.740 ;
        RECT 72.645 95.420 72.965 95.740 ;
        RECT 43.690 89.980 44.010 90.300 ;
        RECT 44.090 89.980 44.410 90.300 ;
        RECT 44.490 89.980 44.810 90.300 ;
        RECT 44.890 89.980 45.210 90.300 ;
        RECT 71.445 89.980 71.765 90.300 ;
        RECT 71.845 89.980 72.165 90.300 ;
        RECT 72.245 89.980 72.565 90.300 ;
        RECT 72.645 89.980 72.965 90.300 ;
        RECT 43.690 84.540 44.010 84.860 ;
        RECT 44.090 84.540 44.410 84.860 ;
        RECT 44.490 84.540 44.810 84.860 ;
        RECT 44.890 84.540 45.210 84.860 ;
        RECT 71.445 84.540 71.765 84.860 ;
        RECT 71.845 84.540 72.165 84.860 ;
        RECT 72.245 84.540 72.565 84.860 ;
        RECT 72.645 84.540 72.965 84.860 ;
        RECT 43.690 79.100 44.010 79.420 ;
        RECT 44.090 79.100 44.410 79.420 ;
        RECT 44.490 79.100 44.810 79.420 ;
        RECT 44.890 79.100 45.210 79.420 ;
        RECT 71.445 79.100 71.765 79.420 ;
        RECT 71.845 79.100 72.165 79.420 ;
        RECT 72.245 79.100 72.565 79.420 ;
        RECT 72.645 79.100 72.965 79.420 ;
        RECT 43.690 73.660 44.010 73.980 ;
        RECT 44.090 73.660 44.410 73.980 ;
        RECT 44.490 73.660 44.810 73.980 ;
        RECT 44.890 73.660 45.210 73.980 ;
        RECT 71.445 73.660 71.765 73.980 ;
        RECT 71.845 73.660 72.165 73.980 ;
        RECT 72.245 73.660 72.565 73.980 ;
        RECT 72.645 73.660 72.965 73.980 ;
        RECT 43.690 68.220 44.010 68.540 ;
        RECT 44.090 68.220 44.410 68.540 ;
        RECT 44.490 68.220 44.810 68.540 ;
        RECT 44.890 68.220 45.210 68.540 ;
        RECT 71.445 68.220 71.765 68.540 ;
        RECT 71.845 68.220 72.165 68.540 ;
        RECT 72.245 68.220 72.565 68.540 ;
        RECT 72.645 68.220 72.965 68.540 ;
        RECT 43.690 62.780 44.010 63.100 ;
        RECT 44.090 62.780 44.410 63.100 ;
        RECT 44.490 62.780 44.810 63.100 ;
        RECT 44.890 62.780 45.210 63.100 ;
        RECT 71.445 62.780 71.765 63.100 ;
        RECT 71.845 62.780 72.165 63.100 ;
        RECT 72.245 62.780 72.565 63.100 ;
        RECT 72.645 62.780 72.965 63.100 ;
        RECT 43.690 57.340 44.010 57.660 ;
        RECT 44.090 57.340 44.410 57.660 ;
        RECT 44.490 57.340 44.810 57.660 ;
        RECT 44.890 57.340 45.210 57.660 ;
        RECT 71.445 57.340 71.765 57.660 ;
        RECT 71.845 57.340 72.165 57.660 ;
        RECT 72.245 57.340 72.565 57.660 ;
        RECT 72.645 57.340 72.965 57.660 ;
        RECT 43.690 51.900 44.010 52.220 ;
        RECT 44.090 51.900 44.410 52.220 ;
        RECT 44.490 51.900 44.810 52.220 ;
        RECT 44.890 51.900 45.210 52.220 ;
        RECT 71.445 51.900 71.765 52.220 ;
        RECT 71.845 51.900 72.165 52.220 ;
        RECT 72.245 51.900 72.565 52.220 ;
        RECT 72.645 51.900 72.965 52.220 ;
        RECT 43.690 46.460 44.010 46.780 ;
        RECT 44.090 46.460 44.410 46.780 ;
        RECT 44.490 46.460 44.810 46.780 ;
        RECT 44.890 46.460 45.210 46.780 ;
        RECT 71.445 46.460 71.765 46.780 ;
        RECT 71.845 46.460 72.165 46.780 ;
        RECT 72.245 46.460 72.565 46.780 ;
        RECT 72.645 46.460 72.965 46.780 ;
        RECT 43.690 41.020 44.010 41.340 ;
        RECT 44.090 41.020 44.410 41.340 ;
        RECT 44.490 41.020 44.810 41.340 ;
        RECT 44.890 41.020 45.210 41.340 ;
        RECT 71.445 41.020 71.765 41.340 ;
        RECT 71.845 41.020 72.165 41.340 ;
        RECT 72.245 41.020 72.565 41.340 ;
        RECT 72.645 41.020 72.965 41.340 ;
        RECT 43.690 35.580 44.010 35.900 ;
        RECT 44.090 35.580 44.410 35.900 ;
        RECT 44.490 35.580 44.810 35.900 ;
        RECT 44.890 35.580 45.210 35.900 ;
        RECT 71.445 35.580 71.765 35.900 ;
        RECT 71.845 35.580 72.165 35.900 ;
        RECT 72.245 35.580 72.565 35.900 ;
        RECT 72.645 35.580 72.965 35.900 ;
        RECT 43.690 30.140 44.010 30.460 ;
        RECT 44.090 30.140 44.410 30.460 ;
        RECT 44.490 30.140 44.810 30.460 ;
        RECT 44.890 30.140 45.210 30.460 ;
        RECT 71.445 30.140 71.765 30.460 ;
        RECT 71.845 30.140 72.165 30.460 ;
        RECT 72.245 30.140 72.565 30.460 ;
        RECT 72.645 30.140 72.965 30.460 ;
        RECT 43.690 24.700 44.010 25.020 ;
        RECT 44.090 24.700 44.410 25.020 ;
        RECT 44.490 24.700 44.810 25.020 ;
        RECT 44.890 24.700 45.210 25.020 ;
        RECT 71.445 24.700 71.765 25.020 ;
        RECT 71.845 24.700 72.165 25.020 ;
        RECT 72.245 24.700 72.565 25.020 ;
        RECT 72.645 24.700 72.965 25.020 ;
        RECT 43.690 19.260 44.010 19.580 ;
        RECT 44.090 19.260 44.410 19.580 ;
        RECT 44.490 19.260 44.810 19.580 ;
        RECT 44.890 19.260 45.210 19.580 ;
        RECT 71.445 19.260 71.765 19.580 ;
        RECT 71.845 19.260 72.165 19.580 ;
        RECT 72.245 19.260 72.565 19.580 ;
        RECT 72.645 19.260 72.965 19.580 ;
      LAYER met4 ;
        RECT 6.600 6.600 8.200 108.400 ;
        RECT 43.650 6.600 45.255 108.400 ;
        RECT 71.405 6.600 73.005 108.400 ;
        RECT 108.460 6.600 110.060 108.400 ;
      LAYER via4 ;
        RECT 6.810 107.010 7.990 108.190 ;
        RECT 6.810 70.270 7.990 71.450 ;
        RECT 6.810 43.070 7.990 44.250 ;
        RECT 6.810 6.810 7.990 7.990 ;
        RECT 43.860 107.010 45.040 108.190 ;
        RECT 43.860 70.270 45.040 71.450 ;
        RECT 43.860 43.070 45.040 44.250 ;
        RECT 43.860 6.810 45.040 7.990 ;
        RECT 71.615 107.010 72.795 108.190 ;
        RECT 71.615 70.270 72.795 71.450 ;
        RECT 71.615 43.070 72.795 44.250 ;
        RECT 71.615 6.810 72.795 7.990 ;
        RECT 108.670 107.010 109.850 108.190 ;
        RECT 108.670 70.270 109.850 71.450 ;
        RECT 108.670 43.070 109.850 44.250 ;
        RECT 108.670 6.810 109.850 7.990 ;
      LAYER met5 ;
        RECT 6.600 106.800 110.060 108.400 ;
        RECT 6.600 70.060 110.060 71.660 ;
        RECT 6.600 42.860 110.060 44.460 ;
        RECT 6.600 6.600 110.060 8.200 ;
    END
  END vssd
  PIN vdda
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3.300 3.300 4.900 111.700 ;
        RECT 33.075 0.000 34.675 115.000 ;
        RECT 60.830 0.000 62.430 115.000 ;
        RECT 88.580 0.000 90.185 115.000 ;
        RECT 111.760 3.300 113.360 111.700 ;
      LAYER via4 ;
        RECT 3.510 110.310 4.690 111.490 ;
        RECT 3.510 87.410 4.690 88.590 ;
        RECT 3.510 60.210 4.690 61.390 ;
        RECT 3.510 33.010 4.690 34.190 ;
        RECT 3.510 3.510 4.690 4.690 ;
        RECT 33.285 110.310 34.465 111.490 ;
        RECT 33.285 87.410 34.465 88.590 ;
        RECT 33.285 60.210 34.465 61.390 ;
        RECT 33.285 33.010 34.465 34.190 ;
        RECT 33.285 3.510 34.465 4.690 ;
        RECT 61.040 110.310 62.220 111.490 ;
        RECT 61.040 87.410 62.220 88.590 ;
        RECT 61.040 60.210 62.220 61.390 ;
        RECT 61.040 33.010 62.220 34.190 ;
        RECT 61.040 3.510 62.220 4.690 ;
        RECT 88.790 110.310 89.970 111.490 ;
        RECT 88.790 87.410 89.970 88.590 ;
        RECT 88.790 60.210 89.970 61.390 ;
        RECT 88.790 33.010 89.970 34.190 ;
        RECT 88.790 3.510 89.970 4.690 ;
        RECT 111.970 110.310 113.150 111.490 ;
        RECT 111.970 87.410 113.150 88.590 ;
        RECT 111.970 60.210 113.150 61.390 ;
        RECT 111.970 33.010 113.150 34.190 ;
        RECT 111.970 3.510 113.150 4.690 ;
      LAYER met5 ;
        RECT 3.300 110.100 113.360 111.700 ;
        RECT 0.000 87.200 116.660 88.800 ;
        RECT 0.000 60.000 116.660 61.600 ;
        RECT 0.000 32.800 116.660 34.400 ;
        RECT 3.300 3.300 113.360 4.900 ;
    END
  END vdda
  PIN vssa
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.600 115.000 ;
        RECT 46.950 0.000 48.555 115.000 ;
        RECT 74.705 0.000 76.305 115.000 ;
        RECT 115.060 0.000 116.660 115.000 ;
      LAYER via4 ;
        RECT 0.210 113.610 1.390 114.790 ;
        RECT 0.210 73.810 1.390 74.990 ;
        RECT 0.210 46.610 1.390 47.790 ;
        RECT 0.210 0.210 1.390 1.390 ;
        RECT 47.160 113.610 48.340 114.790 ;
        RECT 47.160 73.810 48.340 74.990 ;
        RECT 47.160 46.610 48.340 47.790 ;
        RECT 47.160 0.210 48.340 1.390 ;
        RECT 74.915 113.610 76.095 114.790 ;
        RECT 74.915 73.810 76.095 74.990 ;
        RECT 74.915 46.610 76.095 47.790 ;
        RECT 74.915 0.210 76.095 1.390 ;
        RECT 115.270 113.610 116.450 114.790 ;
        RECT 115.270 73.810 116.450 74.990 ;
        RECT 115.270 46.610 116.450 47.790 ;
        RECT 115.270 0.210 116.450 1.390 ;
      LAYER met5 ;
        RECT 0.000 113.400 116.660 115.000 ;
        RECT 0.000 73.600 116.660 75.200 ;
        RECT 0.000 46.400 116.660 48.000 ;
        RECT 0.000 0.000 116.660 1.600 ;
    END
  END vssa
  OBS
      LAYER nwell ;
        RECT 16.510 96.885 100.150 98.490 ;
      LAYER pwell ;
        RECT 31.105 95.900 31.275 96.425 ;
        RECT 45.365 95.900 45.535 96.425 ;
        RECT 59.625 95.900 59.795 96.425 ;
        RECT 73.885 95.900 74.055 96.425 ;
        RECT 88.145 95.900 88.315 96.425 ;
        RECT 16.845 95.495 17.015 95.665 ;
        RECT 18.225 95.495 18.395 95.665 ;
        RECT 19.605 95.495 19.775 95.665 ;
        RECT 20.985 95.495 21.155 95.665 ;
        RECT 23.745 95.495 23.915 95.665 ;
        RECT 26.505 95.495 26.675 95.665 ;
        RECT 29.265 95.495 29.435 95.665 ;
        RECT 30.195 95.520 30.355 95.630 ;
        RECT 31.565 95.495 31.735 95.665 ;
        RECT 32.945 95.495 33.115 95.665 ;
        RECT 37.085 95.495 37.255 95.665 ;
        RECT 38.465 95.495 38.635 95.665 ;
        RECT 42.605 95.495 42.775 95.665 ;
        RECT 43.985 95.495 44.155 95.665 ;
        RECT 45.825 95.495 45.995 95.665 ;
        RECT 49.505 95.495 49.675 95.665 ;
        RECT 51.345 95.495 51.515 95.665 ;
        RECT 55.025 95.495 55.195 95.665 ;
        RECT 56.865 95.495 57.035 95.665 ;
        RECT 58.700 95.525 58.820 95.635 ;
        RECT 59.625 95.495 59.795 95.665 ;
        RECT 60.085 95.495 60.255 95.665 ;
        RECT 61.005 95.495 61.175 95.665 ;
        RECT 65.605 95.495 65.775 95.665 ;
        RECT 66.525 95.495 66.695 95.665 ;
        RECT 71.125 95.495 71.295 95.665 ;
        RECT 72.045 95.495 72.215 95.665 ;
        RECT 74.345 95.495 74.515 95.665 ;
        RECT 77.565 95.495 77.735 95.665 ;
        RECT 79.865 95.495 80.035 95.665 ;
        RECT 83.085 95.495 83.255 95.665 ;
        RECT 85.385 95.495 85.555 95.665 ;
        RECT 86.760 95.525 86.880 95.635 ;
        RECT 87.685 95.495 87.855 95.665 ;
        RECT 88.605 95.495 88.775 95.665 ;
        RECT 89.065 95.495 89.235 95.665 ;
        RECT 92.755 95.520 92.915 95.630 ;
        RECT 93.665 95.495 93.835 95.665 ;
        RECT 94.125 95.495 94.295 95.665 ;
        RECT 95.045 95.495 95.215 95.665 ;
        RECT 97.815 95.530 97.975 95.640 ;
        RECT 99.645 95.495 99.815 95.665 ;
        RECT 31.105 94.735 31.275 95.260 ;
        RECT 59.165 94.735 59.335 95.260 ;
        RECT 87.225 94.735 87.395 95.260 ;
      LAYER nwell ;
        RECT 16.510 91.445 100.150 94.275 ;
      LAYER pwell ;
        RECT 44.905 90.460 45.075 90.985 ;
        RECT 72.965 90.460 73.135 90.985 ;
        RECT 16.845 90.055 17.015 90.225 ;
        RECT 18.225 90.055 18.395 90.225 ;
        RECT 23.745 90.055 23.915 90.225 ;
        RECT 29.265 90.055 29.435 90.225 ;
        RECT 31.565 90.055 31.735 90.225 ;
        RECT 34.785 90.055 34.955 90.225 ;
        RECT 37.085 90.055 37.255 90.225 ;
        RECT 40.305 90.055 40.475 90.225 ;
        RECT 42.605 90.055 42.775 90.225 ;
        RECT 43.995 90.090 44.155 90.200 ;
        RECT 45.365 90.055 45.535 90.225 ;
        RECT 48.125 90.055 48.295 90.225 ;
        RECT 50.885 90.055 51.055 90.225 ;
        RECT 53.645 90.055 53.815 90.225 ;
        RECT 56.405 90.055 56.575 90.225 ;
        RECT 59.625 90.055 59.795 90.225 ;
        RECT 61.925 90.055 62.095 90.225 ;
        RECT 62.385 90.055 62.555 90.225 ;
        RECT 63.760 90.085 63.880 90.195 ;
        RECT 64.225 90.055 64.395 90.225 ;
        RECT 67.445 90.055 67.615 90.225 ;
        RECT 71.125 90.055 71.295 90.225 ;
        RECT 73.425 90.055 73.595 90.225 ;
        RECT 76.645 90.055 76.815 90.225 ;
        RECT 78.945 90.055 79.115 90.225 ;
        RECT 82.165 90.055 82.335 90.225 ;
        RECT 84.465 90.055 84.635 90.225 ;
        RECT 85.845 90.055 86.015 90.225 ;
        RECT 87.685 90.055 87.855 90.225 ;
        RECT 89.985 90.055 90.155 90.225 ;
        RECT 93.205 90.055 93.375 90.225 ;
        RECT 93.665 90.055 93.835 90.225 ;
        RECT 95.045 90.055 95.215 90.225 ;
        RECT 99.645 90.055 99.815 90.225 ;
        RECT 31.105 89.295 31.275 89.820 ;
        RECT 59.165 89.295 59.335 89.820 ;
        RECT 87.225 89.295 87.395 89.820 ;
      LAYER nwell ;
        RECT 16.510 86.005 100.150 88.835 ;
      LAYER pwell ;
        RECT 44.905 85.020 45.075 85.545 ;
        RECT 72.965 85.020 73.135 85.545 ;
        RECT 16.845 84.615 17.015 84.785 ;
        RECT 18.225 84.615 18.395 84.785 ;
        RECT 23.745 84.615 23.915 84.785 ;
        RECT 29.265 84.615 29.435 84.785 ;
        RECT 31.565 84.615 31.735 84.785 ;
        RECT 34.785 84.615 34.955 84.785 ;
        RECT 35.245 84.615 35.415 84.785 ;
        RECT 36.625 84.615 36.795 84.785 ;
        RECT 40.305 84.615 40.475 84.785 ;
        RECT 42.145 84.615 42.315 84.785 ;
        RECT 43.995 84.650 44.155 84.760 ;
        RECT 45.365 84.615 45.535 84.785 ;
        RECT 47.665 84.615 47.835 84.785 ;
        RECT 50.885 84.615 51.055 84.785 ;
        RECT 53.185 84.615 53.355 84.785 ;
        RECT 56.405 84.615 56.575 84.785 ;
        RECT 58.700 84.645 58.820 84.755 ;
        RECT 59.625 84.615 59.795 84.785 ;
        RECT 61.925 84.615 62.095 84.785 ;
        RECT 65.145 84.615 65.315 84.785 ;
        RECT 67.445 84.615 67.615 84.785 ;
        RECT 70.665 84.615 70.835 84.785 ;
        RECT 73.425 84.615 73.595 84.785 ;
        RECT 76.185 84.615 76.355 84.785 ;
        RECT 78.945 84.615 79.115 84.785 ;
        RECT 81.705 84.615 81.875 84.785 ;
        RECT 84.465 84.615 84.635 84.785 ;
        RECT 87.685 84.615 87.855 84.785 ;
        RECT 89.985 84.615 90.155 84.785 ;
        RECT 93.205 84.615 93.375 84.785 ;
        RECT 95.505 84.615 95.675 84.785 ;
        RECT 98.260 84.645 98.380 84.755 ;
        RECT 99.645 84.615 99.815 84.785 ;
        RECT 31.105 83.855 31.275 84.380 ;
        RECT 59.165 83.855 59.335 84.380 ;
        RECT 87.225 83.855 87.395 84.380 ;
      LAYER nwell ;
        RECT 16.510 80.565 100.150 83.395 ;
      LAYER pwell ;
        RECT 44.905 79.580 45.075 80.105 ;
        RECT 72.965 79.580 73.135 80.105 ;
        RECT 16.845 79.175 17.015 79.345 ;
        RECT 18.225 79.175 18.395 79.345 ;
        RECT 23.745 79.175 23.915 79.345 ;
        RECT 29.265 79.175 29.435 79.345 ;
        RECT 31.565 79.175 31.735 79.345 ;
        RECT 34.785 79.175 34.955 79.345 ;
        RECT 37.085 79.175 37.255 79.345 ;
        RECT 37.540 79.205 37.660 79.315 ;
        RECT 38.005 79.175 38.175 79.345 ;
        RECT 38.925 79.175 39.095 79.345 ;
        RECT 41.225 79.175 41.395 79.345 ;
        RECT 45.365 79.175 45.535 79.345 ;
        RECT 47.665 79.175 47.835 79.345 ;
        RECT 50.885 79.175 51.055 79.345 ;
        RECT 53.185 79.175 53.355 79.345 ;
        RECT 56.405 79.175 56.575 79.345 ;
        RECT 58.700 79.205 58.820 79.315 ;
        RECT 59.625 79.175 59.795 79.345 ;
        RECT 61.925 79.175 62.095 79.345 ;
        RECT 65.145 79.175 65.315 79.345 ;
        RECT 67.445 79.175 67.615 79.345 ;
        RECT 70.665 79.175 70.835 79.345 ;
        RECT 73.425 79.175 73.595 79.345 ;
        RECT 78.945 79.175 79.115 79.345 ;
        RECT 82.165 79.175 82.335 79.345 ;
        RECT 84.465 79.175 84.635 79.345 ;
        RECT 85.845 79.175 86.015 79.345 ;
        RECT 87.685 79.175 87.855 79.345 ;
        RECT 89.985 79.175 90.155 79.345 ;
        RECT 93.205 79.175 93.375 79.345 ;
        RECT 95.505 79.175 95.675 79.345 ;
        RECT 98.260 79.205 98.380 79.315 ;
        RECT 99.645 79.175 99.815 79.345 ;
        RECT 31.105 78.415 31.275 78.940 ;
        RECT 59.165 78.415 59.335 78.940 ;
        RECT 87.225 78.415 87.395 78.940 ;
      LAYER nwell ;
        RECT 16.510 75.125 100.150 77.955 ;
      LAYER pwell ;
        RECT 44.905 74.140 45.075 74.665 ;
        RECT 72.965 74.140 73.135 74.665 ;
        RECT 16.845 73.735 17.015 73.905 ;
        RECT 18.225 73.735 18.395 73.905 ;
        RECT 23.745 73.735 23.915 73.905 ;
        RECT 29.265 73.735 29.435 73.905 ;
        RECT 31.565 73.735 31.735 73.905 ;
        RECT 34.785 73.735 34.955 73.905 ;
        RECT 37.085 73.735 37.255 73.905 ;
        RECT 40.305 73.735 40.475 73.905 ;
        RECT 42.605 73.735 42.775 73.905 ;
        RECT 43.995 73.770 44.155 73.880 ;
        RECT 45.365 73.735 45.535 73.905 ;
        RECT 48.125 73.735 48.295 73.905 ;
        RECT 50.885 73.735 51.055 73.905 ;
        RECT 53.645 73.735 53.815 73.905 ;
        RECT 56.405 73.735 56.575 73.905 ;
        RECT 59.625 73.735 59.795 73.905 ;
        RECT 61.925 73.735 62.095 73.905 ;
        RECT 65.145 73.735 65.315 73.905 ;
        RECT 67.445 73.735 67.615 73.905 ;
        RECT 70.665 73.735 70.835 73.905 ;
        RECT 73.425 73.735 73.595 73.905 ;
        RECT 76.185 73.735 76.355 73.905 ;
        RECT 78.945 73.735 79.115 73.905 ;
        RECT 81.705 73.735 81.875 73.905 ;
        RECT 84.465 73.735 84.635 73.905 ;
        RECT 87.685 73.735 87.855 73.905 ;
        RECT 89.985 73.735 90.155 73.905 ;
        RECT 93.205 73.735 93.375 73.905 ;
        RECT 95.505 73.735 95.675 73.905 ;
        RECT 98.260 73.765 98.380 73.875 ;
        RECT 99.645 73.735 99.815 73.905 ;
        RECT 31.105 72.975 31.275 73.500 ;
        RECT 59.165 72.975 59.335 73.500 ;
        RECT 87.225 72.975 87.395 73.500 ;
      LAYER nwell ;
        RECT 16.510 69.685 100.150 72.515 ;
      LAYER pwell ;
        RECT 44.905 68.700 45.075 69.225 ;
        RECT 72.965 68.700 73.135 69.225 ;
        RECT 16.845 68.295 17.015 68.465 ;
        RECT 18.225 68.295 18.395 68.465 ;
        RECT 23.745 68.295 23.915 68.465 ;
        RECT 29.265 68.295 29.435 68.465 ;
        RECT 31.565 68.295 31.735 68.465 ;
        RECT 34.785 68.295 34.955 68.465 ;
        RECT 37.085 68.295 37.255 68.465 ;
        RECT 40.305 68.295 40.475 68.465 ;
        RECT 42.605 68.295 42.775 68.465 ;
        RECT 43.995 68.330 44.155 68.440 ;
        RECT 45.365 68.295 45.535 68.465 ;
        RECT 48.125 68.295 48.295 68.465 ;
        RECT 50.885 68.295 51.055 68.465 ;
        RECT 53.645 68.295 53.815 68.465 ;
        RECT 56.405 68.435 56.575 68.465 ;
        RECT 56.400 68.325 56.575 68.435 ;
        RECT 56.405 68.295 56.575 68.325 ;
        RECT 57.785 68.295 57.955 68.465 ;
        RECT 58.255 68.320 58.415 68.430 ;
        RECT 59.625 68.295 59.795 68.465 ;
        RECT 61.925 68.295 62.095 68.465 ;
        RECT 65.145 68.295 65.315 68.465 ;
        RECT 67.445 68.295 67.615 68.465 ;
        RECT 70.665 68.295 70.835 68.465 ;
        RECT 73.425 68.295 73.595 68.465 ;
        RECT 76.185 68.295 76.355 68.465 ;
        RECT 78.945 68.295 79.115 68.465 ;
        RECT 81.705 68.295 81.875 68.465 ;
        RECT 84.465 68.295 84.635 68.465 ;
        RECT 87.685 68.295 87.855 68.465 ;
        RECT 89.985 68.295 90.155 68.465 ;
        RECT 93.205 68.295 93.375 68.465 ;
        RECT 95.505 68.295 95.675 68.465 ;
        RECT 98.260 68.325 98.380 68.435 ;
        RECT 99.645 68.295 99.815 68.465 ;
        RECT 31.105 67.535 31.275 68.060 ;
        RECT 59.165 67.535 59.335 68.060 ;
        RECT 87.225 67.535 87.395 68.060 ;
      LAYER nwell ;
        RECT 16.510 64.245 100.150 67.075 ;
      LAYER pwell ;
        RECT 44.905 63.260 45.075 63.785 ;
        RECT 72.965 63.260 73.135 63.785 ;
        RECT 16.845 62.855 17.015 63.025 ;
        RECT 18.225 62.855 18.395 63.025 ;
        RECT 19.605 62.855 19.775 63.025 ;
        RECT 20.985 62.855 21.155 63.025 ;
        RECT 23.745 62.855 23.915 63.025 ;
        RECT 26.505 62.855 26.675 63.025 ;
        RECT 29.265 62.855 29.435 63.025 ;
        RECT 30.195 62.880 30.355 62.990 ;
        RECT 31.565 62.855 31.735 63.025 ;
        RECT 34.785 62.855 34.955 63.025 ;
        RECT 37.085 62.855 37.255 63.025 ;
        RECT 40.305 62.855 40.475 63.025 ;
        RECT 40.765 62.855 40.935 63.025 ;
        RECT 43.995 62.890 44.155 63.000 ;
        RECT 45.365 62.855 45.535 63.025 ;
        RECT 49.505 62.855 49.675 63.025 ;
        RECT 50.885 62.855 51.055 63.025 ;
        RECT 55.025 62.855 55.195 63.025 ;
        RECT 56.405 62.855 56.575 63.025 ;
        RECT 60.085 62.995 60.255 63.025 ;
        RECT 58.700 62.885 58.820 62.995 ;
        RECT 59.620 62.885 59.740 62.995 ;
        RECT 60.080 62.885 60.255 62.995 ;
        RECT 60.085 62.855 60.255 62.885 ;
        RECT 60.545 62.855 60.715 63.025 ;
        RECT 61.925 62.855 62.095 63.025 ;
        RECT 67.445 62.855 67.615 63.025 ;
        RECT 68.825 62.855 68.995 63.025 ;
        RECT 69.285 62.855 69.455 63.025 ;
        RECT 73.425 62.855 73.595 63.025 ;
        RECT 77.565 62.855 77.735 63.025 ;
        RECT 78.945 62.855 79.115 63.025 ;
        RECT 83.085 62.855 83.255 63.025 ;
        RECT 84.465 62.855 84.635 63.025 ;
        RECT 86.760 62.885 86.880 62.995 ;
        RECT 87.685 62.855 87.855 63.025 ;
        RECT 89.985 62.855 90.155 63.025 ;
        RECT 93.205 62.855 93.375 63.025 ;
        RECT 95.505 62.855 95.675 63.025 ;
        RECT 98.260 62.885 98.380 62.995 ;
        RECT 99.645 62.855 99.815 63.025 ;
        RECT 31.105 62.095 31.275 62.620 ;
        RECT 59.165 62.095 59.335 62.620 ;
        RECT 87.225 62.095 87.395 62.620 ;
      LAYER nwell ;
        RECT 16.510 58.805 100.150 61.635 ;
      LAYER pwell ;
        RECT 44.905 57.820 45.075 58.345 ;
        RECT 72.965 57.820 73.135 58.345 ;
        RECT 16.845 57.415 17.015 57.585 ;
        RECT 18.225 57.415 18.395 57.585 ;
        RECT 23.745 57.415 23.915 57.585 ;
        RECT 29.265 57.415 29.435 57.585 ;
        RECT 31.565 57.415 31.735 57.585 ;
        RECT 34.785 57.415 34.955 57.585 ;
        RECT 37.085 57.415 37.255 57.585 ;
        RECT 37.540 57.445 37.660 57.555 ;
        RECT 38.005 57.415 38.175 57.585 ;
        RECT 41.225 57.415 41.395 57.585 ;
        RECT 42.605 57.415 42.775 57.585 ;
        RECT 45.365 57.415 45.535 57.585 ;
        RECT 48.125 57.415 48.295 57.585 ;
        RECT 50.885 57.415 51.055 57.585 ;
        RECT 53.645 57.415 53.815 57.585 ;
        RECT 56.405 57.415 56.575 57.585 ;
        RECT 59.625 57.415 59.795 57.585 ;
        RECT 61.925 57.415 62.095 57.585 ;
        RECT 63.765 57.415 63.935 57.585 ;
        RECT 65.145 57.415 65.315 57.585 ;
        RECT 66.985 57.415 67.155 57.585 ;
        RECT 68.365 57.415 68.535 57.585 ;
        RECT 72.500 57.445 72.620 57.555 ;
        RECT 73.425 57.415 73.595 57.585 ;
        RECT 73.885 57.415 74.055 57.585 ;
        RECT 78.945 57.415 79.115 57.585 ;
        RECT 79.405 57.415 79.575 57.585 ;
        RECT 84.465 57.415 84.635 57.585 ;
        RECT 84.925 57.415 85.095 57.585 ;
        RECT 86.760 57.445 86.880 57.555 ;
        RECT 87.685 57.415 87.855 57.585 ;
        RECT 89.985 57.415 90.155 57.585 ;
        RECT 93.205 57.415 93.375 57.585 ;
        RECT 95.505 57.415 95.675 57.585 ;
        RECT 98.260 57.445 98.380 57.555 ;
        RECT 99.645 57.415 99.815 57.585 ;
        RECT 31.105 56.655 31.275 57.180 ;
        RECT 59.165 56.655 59.335 57.180 ;
        RECT 87.225 56.655 87.395 57.180 ;
      LAYER nwell ;
        RECT 16.510 53.365 100.150 56.195 ;
      LAYER pwell ;
        RECT 44.905 52.380 45.075 52.905 ;
        RECT 72.965 52.380 73.135 52.905 ;
        RECT 16.845 51.975 17.015 52.145 ;
        RECT 18.225 51.975 18.395 52.145 ;
        RECT 23.745 51.975 23.915 52.145 ;
        RECT 29.265 51.975 29.435 52.145 ;
        RECT 31.565 51.975 31.735 52.145 ;
        RECT 34.785 51.975 34.955 52.145 ;
        RECT 37.085 51.975 37.255 52.145 ;
        RECT 40.305 51.975 40.475 52.145 ;
        RECT 42.605 51.975 42.775 52.145 ;
        RECT 43.995 52.010 44.155 52.120 ;
        RECT 45.365 51.975 45.535 52.145 ;
        RECT 48.125 51.975 48.295 52.145 ;
        RECT 50.885 51.975 51.055 52.145 ;
        RECT 53.645 51.975 53.815 52.145 ;
        RECT 56.405 51.975 56.575 52.145 ;
        RECT 59.625 51.975 59.795 52.145 ;
        RECT 61.005 51.975 61.175 52.145 ;
        RECT 65.605 51.975 65.775 52.145 ;
        RECT 69.745 51.975 69.915 52.145 ;
        RECT 71.125 51.975 71.295 52.145 ;
        RECT 73.425 51.975 73.595 52.145 ;
        RECT 75.265 51.975 75.435 52.145 ;
        RECT 78.945 51.975 79.115 52.145 ;
        RECT 80.785 51.975 80.955 52.145 ;
        RECT 84.465 51.975 84.635 52.145 ;
        RECT 86.315 52.000 86.475 52.110 ;
        RECT 87.685 51.975 87.855 52.145 ;
        RECT 89.985 51.975 90.155 52.145 ;
        RECT 93.205 51.975 93.375 52.145 ;
        RECT 95.505 51.975 95.675 52.145 ;
        RECT 98.260 52.005 98.380 52.115 ;
        RECT 99.645 51.975 99.815 52.145 ;
        RECT 31.105 51.215 31.275 51.740 ;
        RECT 59.165 51.215 59.335 51.740 ;
        RECT 87.225 51.215 87.395 51.740 ;
      LAYER nwell ;
        RECT 16.510 47.925 100.150 50.755 ;
      LAYER pwell ;
        RECT 44.905 46.940 45.075 47.465 ;
        RECT 72.965 46.940 73.135 47.465 ;
        RECT 16.845 46.535 17.015 46.705 ;
        RECT 18.225 46.535 18.395 46.705 ;
        RECT 19.605 46.535 19.775 46.705 ;
        RECT 20.985 46.535 21.155 46.705 ;
        RECT 23.745 46.535 23.915 46.705 ;
        RECT 26.505 46.535 26.675 46.705 ;
        RECT 29.265 46.535 29.435 46.705 ;
        RECT 31.565 46.535 31.735 46.705 ;
        RECT 32.025 46.535 32.195 46.705 ;
        RECT 37.085 46.535 37.255 46.705 ;
        RECT 37.545 46.535 37.715 46.705 ;
        RECT 42.605 46.535 42.775 46.705 ;
        RECT 43.065 46.535 43.235 46.705 ;
        RECT 45.365 46.535 45.535 46.705 ;
        RECT 48.125 46.535 48.295 46.705 ;
        RECT 50.885 46.535 51.055 46.705 ;
        RECT 53.645 46.535 53.815 46.705 ;
        RECT 56.405 46.535 56.575 46.705 ;
        RECT 59.160 46.565 59.280 46.675 ;
        RECT 59.625 46.535 59.795 46.705 ;
        RECT 60.545 46.535 60.715 46.705 ;
        RECT 61.005 46.535 61.175 46.705 ;
        RECT 62.845 46.535 63.015 46.705 ;
        RECT 66.525 46.535 66.695 46.705 ;
        RECT 68.365 46.535 68.535 46.705 ;
        RECT 72.055 46.570 72.215 46.680 ;
        RECT 73.425 46.535 73.595 46.705 ;
        RECT 73.885 46.535 74.055 46.705 ;
        RECT 78.945 46.535 79.115 46.705 ;
        RECT 79.405 46.535 79.575 46.705 ;
        RECT 84.465 46.535 84.635 46.705 ;
        RECT 84.925 46.535 85.095 46.705 ;
        RECT 86.760 46.565 86.880 46.675 ;
        RECT 87.685 46.535 87.855 46.705 ;
        RECT 89.985 46.535 90.155 46.705 ;
        RECT 93.205 46.535 93.375 46.705 ;
        RECT 95.505 46.535 95.675 46.705 ;
        RECT 98.260 46.565 98.380 46.675 ;
        RECT 99.645 46.535 99.815 46.705 ;
        RECT 31.105 45.775 31.275 46.300 ;
        RECT 59.165 45.775 59.335 46.300 ;
        RECT 87.225 45.775 87.395 46.300 ;
      LAYER nwell ;
        RECT 16.510 42.485 100.150 45.315 ;
      LAYER pwell ;
        RECT 44.905 41.500 45.075 42.025 ;
        RECT 72.965 41.500 73.135 42.025 ;
        RECT 16.845 41.095 17.015 41.265 ;
        RECT 18.225 41.095 18.395 41.265 ;
        RECT 23.745 41.095 23.915 41.265 ;
        RECT 29.265 41.095 29.435 41.265 ;
        RECT 31.565 41.095 31.735 41.265 ;
        RECT 34.785 41.095 34.955 41.265 ;
        RECT 37.085 41.095 37.255 41.265 ;
        RECT 40.305 41.095 40.475 41.265 ;
        RECT 42.605 41.095 42.775 41.265 ;
        RECT 43.995 41.130 44.155 41.240 ;
        RECT 45.365 41.095 45.535 41.265 ;
        RECT 48.125 41.095 48.295 41.265 ;
        RECT 50.885 41.095 51.055 41.265 ;
        RECT 53.645 41.095 53.815 41.265 ;
        RECT 56.405 41.095 56.575 41.265 ;
        RECT 59.625 41.095 59.795 41.265 ;
        RECT 61.925 41.095 62.095 41.265 ;
        RECT 65.145 41.095 65.315 41.265 ;
        RECT 67.445 41.095 67.615 41.265 ;
        RECT 70.665 41.095 70.835 41.265 ;
        RECT 73.425 41.095 73.595 41.265 ;
        RECT 76.185 41.095 76.355 41.265 ;
        RECT 78.945 41.095 79.115 41.265 ;
        RECT 81.705 41.095 81.875 41.265 ;
        RECT 84.465 41.095 84.635 41.265 ;
        RECT 87.685 41.095 87.855 41.265 ;
        RECT 89.985 41.095 90.155 41.265 ;
        RECT 93.205 41.095 93.375 41.265 ;
        RECT 95.505 41.095 95.675 41.265 ;
        RECT 98.260 41.125 98.380 41.235 ;
        RECT 99.645 41.095 99.815 41.265 ;
        RECT 31.105 40.335 31.275 40.860 ;
        RECT 59.165 40.335 59.335 40.860 ;
        RECT 87.225 40.335 87.395 40.860 ;
      LAYER nwell ;
        RECT 16.510 37.045 100.150 39.875 ;
      LAYER pwell ;
        RECT 44.905 36.060 45.075 36.585 ;
        RECT 72.965 36.060 73.135 36.585 ;
        RECT 16.845 35.655 17.015 35.825 ;
        RECT 18.225 35.655 18.395 35.825 ;
        RECT 19.605 35.655 19.775 35.825 ;
        RECT 20.985 35.655 21.155 35.825 ;
        RECT 23.745 35.655 23.915 35.825 ;
        RECT 26.505 35.655 26.675 35.825 ;
        RECT 29.265 35.655 29.435 35.825 ;
        RECT 30.195 35.680 30.355 35.790 ;
        RECT 31.565 35.655 31.735 35.825 ;
        RECT 34.785 35.655 34.955 35.825 ;
        RECT 37.085 35.655 37.255 35.825 ;
        RECT 40.305 35.655 40.475 35.825 ;
        RECT 42.605 35.655 42.775 35.825 ;
        RECT 43.995 35.690 44.155 35.800 ;
        RECT 45.365 35.655 45.535 35.825 ;
        RECT 48.125 35.655 48.295 35.825 ;
        RECT 50.885 35.655 51.055 35.825 ;
        RECT 53.645 35.655 53.815 35.825 ;
        RECT 56.405 35.655 56.575 35.825 ;
        RECT 59.625 35.655 59.795 35.825 ;
        RECT 61.925 35.655 62.095 35.825 ;
        RECT 65.145 35.655 65.315 35.825 ;
        RECT 67.445 35.655 67.615 35.825 ;
        RECT 70.665 35.655 70.835 35.825 ;
        RECT 73.425 35.655 73.595 35.825 ;
        RECT 76.185 35.655 76.355 35.825 ;
        RECT 78.945 35.655 79.115 35.825 ;
        RECT 81.705 35.655 81.875 35.825 ;
        RECT 84.465 35.655 84.635 35.825 ;
        RECT 87.685 35.655 87.855 35.825 ;
        RECT 89.985 35.655 90.155 35.825 ;
        RECT 93.205 35.655 93.375 35.825 ;
        RECT 93.665 35.655 93.835 35.825 ;
        RECT 95.045 35.655 95.215 35.825 ;
        RECT 99.645 35.655 99.815 35.825 ;
        RECT 31.105 34.895 31.275 35.420 ;
        RECT 59.165 34.895 59.335 35.420 ;
        RECT 87.225 34.895 87.395 35.420 ;
      LAYER nwell ;
        RECT 16.510 31.605 100.150 34.435 ;
      LAYER pwell ;
        RECT 44.905 30.620 45.075 31.145 ;
        RECT 72.965 30.620 73.135 31.145 ;
        RECT 16.845 30.215 17.015 30.385 ;
        RECT 18.225 30.215 18.395 30.385 ;
        RECT 23.745 30.215 23.915 30.385 ;
        RECT 29.265 30.215 29.435 30.385 ;
        RECT 31.565 30.215 31.735 30.385 ;
        RECT 34.785 30.215 34.955 30.385 ;
        RECT 37.085 30.215 37.255 30.385 ;
        RECT 40.305 30.215 40.475 30.385 ;
        RECT 42.605 30.215 42.775 30.385 ;
        RECT 43.995 30.250 44.155 30.360 ;
        RECT 45.365 30.215 45.535 30.385 ;
        RECT 48.125 30.215 48.295 30.385 ;
        RECT 50.885 30.215 51.055 30.385 ;
        RECT 53.645 30.215 53.815 30.385 ;
        RECT 56.405 30.215 56.575 30.385 ;
        RECT 59.625 30.215 59.795 30.385 ;
        RECT 61.925 30.215 62.095 30.385 ;
        RECT 65.145 30.215 65.315 30.385 ;
        RECT 67.445 30.215 67.615 30.385 ;
        RECT 70.665 30.215 70.835 30.385 ;
        RECT 73.425 30.215 73.595 30.385 ;
        RECT 76.185 30.215 76.355 30.385 ;
        RECT 78.945 30.215 79.115 30.385 ;
        RECT 81.705 30.215 81.875 30.385 ;
        RECT 84.465 30.215 84.635 30.385 ;
        RECT 87.685 30.215 87.855 30.385 ;
        RECT 89.985 30.215 90.155 30.385 ;
        RECT 93.205 30.215 93.375 30.385 ;
        RECT 95.505 30.215 95.675 30.385 ;
        RECT 98.260 30.245 98.380 30.355 ;
        RECT 99.645 30.215 99.815 30.385 ;
        RECT 31.105 29.455 31.275 29.980 ;
        RECT 59.165 29.455 59.335 29.980 ;
        RECT 87.225 29.455 87.395 29.980 ;
      LAYER nwell ;
        RECT 16.510 26.165 100.150 28.995 ;
      LAYER pwell ;
        RECT 44.905 25.180 45.075 25.705 ;
        RECT 72.965 25.180 73.135 25.705 ;
        RECT 16.845 24.775 17.015 24.945 ;
        RECT 18.225 24.775 18.395 24.945 ;
        RECT 23.745 24.775 23.915 24.945 ;
        RECT 29.265 24.775 29.435 24.945 ;
        RECT 31.565 24.775 31.735 24.945 ;
        RECT 34.785 24.775 34.955 24.945 ;
        RECT 37.085 24.775 37.255 24.945 ;
        RECT 40.305 24.775 40.475 24.945 ;
        RECT 42.605 24.775 42.775 24.945 ;
        RECT 43.995 24.810 44.155 24.920 ;
        RECT 45.365 24.775 45.535 24.945 ;
        RECT 48.125 24.775 48.295 24.945 ;
        RECT 50.885 24.775 51.055 24.945 ;
        RECT 53.645 24.775 53.815 24.945 ;
        RECT 56.405 24.775 56.575 24.945 ;
        RECT 59.625 24.775 59.795 24.945 ;
        RECT 61.925 24.775 62.095 24.945 ;
        RECT 65.145 24.775 65.315 24.945 ;
        RECT 67.445 24.775 67.615 24.945 ;
        RECT 70.665 24.775 70.835 24.945 ;
        RECT 72.500 24.805 72.620 24.915 ;
        RECT 72.965 24.775 73.135 24.945 ;
        RECT 73.425 24.775 73.595 24.945 ;
        RECT 76.185 24.775 76.355 24.945 ;
        RECT 78.945 24.775 79.115 24.945 ;
        RECT 81.705 24.775 81.875 24.945 ;
        RECT 84.465 24.775 84.635 24.945 ;
        RECT 87.685 24.775 87.855 24.945 ;
        RECT 89.985 24.775 90.155 24.945 ;
        RECT 93.205 24.775 93.375 24.945 ;
        RECT 95.505 24.775 95.675 24.945 ;
        RECT 98.260 24.805 98.380 24.915 ;
        RECT 99.645 24.775 99.815 24.945 ;
        RECT 31.105 24.015 31.275 24.540 ;
        RECT 59.165 24.015 59.335 24.540 ;
        RECT 87.225 24.015 87.395 24.540 ;
      LAYER nwell ;
        RECT 16.510 20.725 100.150 23.555 ;
      LAYER pwell ;
        RECT 44.905 19.740 45.075 20.265 ;
        RECT 72.965 19.740 73.135 20.265 ;
        RECT 16.845 19.335 17.015 19.505 ;
        RECT 18.225 19.335 18.395 19.505 ;
        RECT 19.605 19.335 19.775 19.505 ;
        RECT 20.985 19.335 21.155 19.505 ;
        RECT 23.745 19.335 23.915 19.505 ;
        RECT 26.505 19.335 26.675 19.505 ;
        RECT 29.265 19.335 29.435 19.505 ;
        RECT 31.565 19.335 31.735 19.505 ;
        RECT 32.025 19.335 32.195 19.505 ;
        RECT 32.945 19.335 33.115 19.505 ;
        RECT 37.545 19.335 37.715 19.505 ;
        RECT 38.465 19.335 38.635 19.505 ;
        RECT 43.065 19.335 43.235 19.505 ;
        RECT 43.985 19.335 44.155 19.505 ;
        RECT 45.365 19.335 45.535 19.505 ;
        RECT 45.825 19.335 45.995 19.505 ;
        RECT 48.580 19.365 48.700 19.475 ;
        RECT 49.045 19.335 49.215 19.505 ;
        RECT 50.425 19.335 50.595 19.505 ;
        RECT 50.885 19.335 51.055 19.505 ;
        RECT 53.640 19.365 53.760 19.475 ;
        RECT 54.105 19.335 54.275 19.505 ;
        RECT 55.945 19.335 56.115 19.505 ;
        RECT 60.085 19.335 60.255 19.505 ;
        RECT 62.845 19.335 63.015 19.505 ;
        RECT 63.305 19.335 63.475 19.505 ;
        RECT 68.365 19.335 68.535 19.505 ;
        RECT 68.825 19.335 68.995 19.505 ;
        RECT 72.055 19.370 72.215 19.480 ;
        RECT 72.505 19.335 72.675 19.505 ;
        RECT 73.425 19.335 73.595 19.505 ;
        RECT 74.345 19.335 74.515 19.505 ;
        RECT 79.865 19.335 80.035 19.505 ;
        RECT 82.165 19.335 82.335 19.505 ;
        RECT 85.385 19.335 85.555 19.505 ;
        RECT 87.685 19.335 87.855 19.505 ;
        RECT 88.605 19.335 88.775 19.505 ;
        RECT 89.985 19.335 90.155 19.505 ;
        RECT 93.205 19.335 93.375 19.505 ;
        RECT 93.665 19.335 93.835 19.505 ;
        RECT 95.045 19.335 95.215 19.505 ;
        RECT 99.645 19.335 99.815 19.505 ;
        RECT 31.105 18.575 31.275 19.100 ;
        RECT 45.365 18.575 45.535 19.100 ;
        RECT 59.625 18.575 59.795 19.100 ;
        RECT 73.885 18.575 74.055 19.100 ;
        RECT 88.145 18.575 88.315 19.100 ;
      LAYER nwell ;
        RECT 16.510 16.510 100.150 18.115 ;
      LAYER li1 ;
        RECT 16.700 98.215 16.845 98.385 ;
        RECT 17.015 98.215 17.305 98.385 ;
        RECT 17.475 98.215 17.765 98.385 ;
        RECT 17.935 98.215 18.225 98.385 ;
        RECT 18.395 98.215 18.685 98.385 ;
        RECT 18.855 98.215 19.145 98.385 ;
        RECT 19.315 98.215 19.605 98.385 ;
        RECT 19.775 98.215 20.065 98.385 ;
        RECT 20.235 98.215 20.525 98.385 ;
        RECT 20.695 98.215 20.985 98.385 ;
        RECT 21.155 98.215 21.445 98.385 ;
        RECT 21.615 98.215 21.905 98.385 ;
        RECT 22.075 98.215 22.365 98.385 ;
        RECT 22.535 98.215 22.825 98.385 ;
        RECT 22.995 98.215 23.285 98.385 ;
        RECT 23.455 98.215 23.745 98.385 ;
        RECT 23.915 98.215 24.205 98.385 ;
        RECT 24.375 98.215 24.665 98.385 ;
        RECT 24.835 98.215 25.125 98.385 ;
        RECT 25.295 98.215 25.585 98.385 ;
        RECT 25.755 98.215 26.045 98.385 ;
        RECT 26.215 98.215 26.505 98.385 ;
        RECT 26.675 98.215 26.965 98.385 ;
        RECT 27.135 98.215 27.425 98.385 ;
        RECT 27.595 98.215 27.885 98.385 ;
        RECT 28.055 98.215 28.345 98.385 ;
        RECT 28.515 98.215 28.805 98.385 ;
        RECT 28.975 98.215 29.265 98.385 ;
        RECT 29.435 98.215 29.725 98.385 ;
        RECT 29.895 98.215 30.185 98.385 ;
        RECT 30.355 98.215 30.645 98.385 ;
        RECT 30.815 98.215 31.105 98.385 ;
        RECT 31.275 98.215 31.565 98.385 ;
        RECT 31.735 98.215 32.025 98.385 ;
        RECT 32.195 98.215 32.485 98.385 ;
        RECT 32.655 98.215 32.945 98.385 ;
        RECT 33.115 98.215 33.405 98.385 ;
        RECT 33.575 98.215 33.865 98.385 ;
        RECT 34.035 98.215 34.325 98.385 ;
        RECT 34.495 98.215 34.785 98.385 ;
        RECT 34.955 98.215 35.245 98.385 ;
        RECT 35.415 98.215 35.705 98.385 ;
        RECT 35.875 98.215 36.165 98.385 ;
        RECT 36.335 98.215 36.625 98.385 ;
        RECT 36.795 98.215 37.085 98.385 ;
        RECT 37.255 98.215 37.545 98.385 ;
        RECT 37.715 98.215 38.005 98.385 ;
        RECT 38.175 98.215 38.465 98.385 ;
        RECT 38.635 98.215 38.925 98.385 ;
        RECT 39.095 98.215 39.385 98.385 ;
        RECT 39.555 98.215 39.845 98.385 ;
        RECT 40.015 98.215 40.305 98.385 ;
        RECT 40.475 98.215 40.765 98.385 ;
        RECT 40.935 98.215 41.225 98.385 ;
        RECT 41.395 98.215 41.685 98.385 ;
        RECT 41.855 98.215 42.145 98.385 ;
        RECT 42.315 98.215 42.605 98.385 ;
        RECT 42.775 98.215 43.065 98.385 ;
        RECT 43.235 98.215 43.525 98.385 ;
        RECT 43.695 98.215 43.985 98.385 ;
        RECT 44.155 98.215 44.445 98.385 ;
        RECT 44.615 98.215 44.905 98.385 ;
        RECT 45.075 98.215 45.365 98.385 ;
        RECT 45.535 98.215 45.825 98.385 ;
        RECT 45.995 98.215 46.285 98.385 ;
        RECT 46.455 98.215 46.745 98.385 ;
        RECT 46.915 98.215 47.205 98.385 ;
        RECT 47.375 98.215 47.665 98.385 ;
        RECT 47.835 98.215 48.125 98.385 ;
        RECT 48.295 98.215 48.585 98.385 ;
        RECT 48.755 98.215 49.045 98.385 ;
        RECT 49.215 98.215 49.505 98.385 ;
        RECT 49.675 98.215 49.965 98.385 ;
        RECT 50.135 98.215 50.425 98.385 ;
        RECT 50.595 98.215 50.885 98.385 ;
        RECT 51.055 98.215 51.345 98.385 ;
        RECT 51.515 98.215 51.805 98.385 ;
        RECT 51.975 98.215 52.265 98.385 ;
        RECT 52.435 98.215 52.725 98.385 ;
        RECT 52.895 98.215 53.185 98.385 ;
        RECT 53.355 98.215 53.645 98.385 ;
        RECT 53.815 98.215 54.105 98.385 ;
        RECT 54.275 98.215 54.565 98.385 ;
        RECT 54.735 98.215 55.025 98.385 ;
        RECT 55.195 98.215 55.485 98.385 ;
        RECT 55.655 98.215 55.945 98.385 ;
        RECT 56.115 98.215 56.405 98.385 ;
        RECT 56.575 98.215 56.865 98.385 ;
        RECT 57.035 98.215 57.325 98.385 ;
        RECT 57.495 98.215 57.785 98.385 ;
        RECT 57.955 98.215 58.245 98.385 ;
        RECT 58.415 98.215 58.705 98.385 ;
        RECT 58.875 98.215 59.165 98.385 ;
        RECT 59.335 98.215 59.625 98.385 ;
        RECT 59.795 98.215 60.085 98.385 ;
        RECT 60.255 98.215 60.545 98.385 ;
        RECT 60.715 98.215 61.005 98.385 ;
        RECT 61.175 98.215 61.465 98.385 ;
        RECT 61.635 98.215 61.925 98.385 ;
        RECT 62.095 98.215 62.385 98.385 ;
        RECT 62.555 98.215 62.845 98.385 ;
        RECT 63.015 98.215 63.305 98.385 ;
        RECT 63.475 98.215 63.765 98.385 ;
        RECT 63.935 98.215 64.225 98.385 ;
        RECT 64.395 98.215 64.685 98.385 ;
        RECT 64.855 98.215 65.145 98.385 ;
        RECT 65.315 98.215 65.605 98.385 ;
        RECT 65.775 98.215 66.065 98.385 ;
        RECT 66.235 98.215 66.525 98.385 ;
        RECT 66.695 98.215 66.985 98.385 ;
        RECT 67.155 98.215 67.445 98.385 ;
        RECT 67.615 98.215 67.905 98.385 ;
        RECT 68.075 98.215 68.365 98.385 ;
        RECT 68.535 98.215 68.825 98.385 ;
        RECT 68.995 98.215 69.285 98.385 ;
        RECT 69.455 98.215 69.745 98.385 ;
        RECT 69.915 98.215 70.205 98.385 ;
        RECT 70.375 98.215 70.665 98.385 ;
        RECT 70.835 98.215 71.125 98.385 ;
        RECT 71.295 98.215 71.585 98.385 ;
        RECT 71.755 98.215 72.045 98.385 ;
        RECT 72.215 98.215 72.505 98.385 ;
        RECT 72.675 98.215 72.965 98.385 ;
        RECT 73.135 98.215 73.425 98.385 ;
        RECT 73.595 98.215 73.885 98.385 ;
        RECT 74.055 98.215 74.345 98.385 ;
        RECT 74.515 98.215 74.805 98.385 ;
        RECT 74.975 98.215 75.265 98.385 ;
        RECT 75.435 98.215 75.725 98.385 ;
        RECT 75.895 98.215 76.185 98.385 ;
        RECT 76.355 98.215 76.645 98.385 ;
        RECT 76.815 98.215 77.105 98.385 ;
        RECT 77.275 98.215 77.565 98.385 ;
        RECT 77.735 98.215 78.025 98.385 ;
        RECT 78.195 98.215 78.485 98.385 ;
        RECT 78.655 98.215 78.945 98.385 ;
        RECT 79.115 98.215 79.405 98.385 ;
        RECT 79.575 98.215 79.865 98.385 ;
        RECT 80.035 98.215 80.325 98.385 ;
        RECT 80.495 98.215 80.785 98.385 ;
        RECT 80.955 98.215 81.245 98.385 ;
        RECT 81.415 98.215 81.705 98.385 ;
        RECT 81.875 98.215 82.165 98.385 ;
        RECT 82.335 98.215 82.625 98.385 ;
        RECT 82.795 98.215 83.085 98.385 ;
        RECT 83.255 98.215 83.545 98.385 ;
        RECT 83.715 98.215 84.005 98.385 ;
        RECT 84.175 98.215 84.465 98.385 ;
        RECT 84.635 98.215 84.925 98.385 ;
        RECT 85.095 98.215 85.385 98.385 ;
        RECT 85.555 98.215 85.845 98.385 ;
        RECT 86.015 98.215 86.305 98.385 ;
        RECT 86.475 98.215 86.765 98.385 ;
        RECT 86.935 98.215 87.225 98.385 ;
        RECT 87.395 98.215 87.685 98.385 ;
        RECT 87.855 98.215 88.145 98.385 ;
        RECT 88.315 98.215 88.605 98.385 ;
        RECT 88.775 98.215 89.065 98.385 ;
        RECT 89.235 98.215 89.525 98.385 ;
        RECT 89.695 98.215 89.985 98.385 ;
        RECT 90.155 98.215 90.445 98.385 ;
        RECT 90.615 98.215 90.905 98.385 ;
        RECT 91.075 98.215 91.365 98.385 ;
        RECT 91.535 98.215 91.825 98.385 ;
        RECT 91.995 98.215 92.285 98.385 ;
        RECT 92.455 98.215 92.745 98.385 ;
        RECT 92.915 98.215 93.205 98.385 ;
        RECT 93.375 98.215 93.665 98.385 ;
        RECT 93.835 98.215 94.125 98.385 ;
        RECT 94.295 98.215 94.585 98.385 ;
        RECT 94.755 98.215 95.045 98.385 ;
        RECT 95.215 98.215 95.505 98.385 ;
        RECT 95.675 98.215 95.965 98.385 ;
        RECT 96.135 98.215 96.425 98.385 ;
        RECT 96.595 98.215 96.885 98.385 ;
        RECT 97.055 98.215 97.345 98.385 ;
        RECT 97.515 98.215 97.805 98.385 ;
        RECT 97.975 98.215 98.265 98.385 ;
        RECT 98.435 98.215 98.725 98.385 ;
        RECT 98.895 98.215 99.185 98.385 ;
        RECT 99.355 98.215 99.645 98.385 ;
        RECT 99.815 98.215 99.960 98.385 ;
        RECT 16.785 97.125 17.995 98.215 ;
        RECT 18.165 97.125 23.510 98.215 ;
        RECT 23.685 97.125 29.030 98.215 ;
        RECT 29.205 97.125 30.875 98.215 ;
        RECT 16.785 96.415 17.305 96.955 ;
        RECT 17.475 96.585 17.995 97.125 ;
        RECT 18.165 96.435 20.745 96.955 ;
        RECT 20.915 96.605 23.510 97.125 ;
        RECT 23.685 96.435 26.265 96.955 ;
        RECT 26.435 96.605 29.030 97.125 ;
        RECT 29.205 96.435 29.955 96.955 ;
        RECT 30.125 96.605 30.875 97.125 ;
        RECT 31.045 97.050 31.335 98.215 ;
        RECT 31.505 97.125 36.850 98.215 ;
        RECT 37.025 97.125 42.370 98.215 ;
        RECT 42.545 97.125 45.135 98.215 ;
        RECT 31.505 96.435 34.085 96.955 ;
        RECT 34.255 96.605 36.850 97.125 ;
        RECT 37.025 96.435 39.605 96.955 ;
        RECT 39.775 96.605 42.370 97.125 ;
        RECT 42.545 96.435 43.755 96.955 ;
        RECT 43.925 96.605 45.135 97.125 ;
        RECT 45.305 97.050 45.595 98.215 ;
        RECT 45.765 97.125 51.110 98.215 ;
        RECT 51.285 97.125 56.630 98.215 ;
        RECT 56.805 97.125 59.395 98.215 ;
        RECT 45.765 96.435 48.345 96.955 ;
        RECT 48.515 96.605 51.110 97.125 ;
        RECT 51.285 96.435 53.865 96.955 ;
        RECT 54.035 96.605 56.630 97.125 ;
        RECT 56.805 96.435 58.015 96.955 ;
        RECT 58.185 96.605 59.395 97.125 ;
        RECT 59.565 97.050 59.855 98.215 ;
        RECT 60.025 97.125 65.370 98.215 ;
        RECT 65.545 97.125 70.890 98.215 ;
        RECT 71.065 97.125 73.655 98.215 ;
        RECT 60.025 96.435 62.605 96.955 ;
        RECT 62.775 96.605 65.370 97.125 ;
        RECT 65.545 96.435 68.125 96.955 ;
        RECT 68.295 96.605 70.890 97.125 ;
        RECT 71.065 96.435 72.275 96.955 ;
        RECT 72.445 96.605 73.655 97.125 ;
        RECT 73.825 97.050 74.115 98.215 ;
        RECT 74.285 97.125 79.630 98.215 ;
        RECT 79.805 97.125 85.150 98.215 ;
        RECT 85.325 97.125 87.915 98.215 ;
        RECT 74.285 96.435 76.865 96.955 ;
        RECT 77.035 96.605 79.630 97.125 ;
        RECT 79.805 96.435 82.385 96.955 ;
        RECT 82.555 96.605 85.150 97.125 ;
        RECT 85.325 96.435 86.535 96.955 ;
        RECT 86.705 96.605 87.915 97.125 ;
        RECT 88.085 97.050 88.375 98.215 ;
        RECT 88.545 97.125 93.890 98.215 ;
        RECT 94.065 97.125 97.575 98.215 ;
        RECT 88.545 96.435 91.125 96.955 ;
        RECT 91.295 96.605 93.890 97.125 ;
        RECT 94.065 96.435 95.715 96.955 ;
        RECT 95.885 96.605 97.575 97.125 ;
        RECT 98.665 97.125 99.875 98.215 ;
        RECT 98.665 96.585 99.185 97.125 ;
        RECT 16.785 95.665 17.995 96.415 ;
        RECT 18.165 95.665 23.510 96.435 ;
        RECT 23.685 95.665 29.030 96.435 ;
        RECT 29.205 95.665 30.875 96.435 ;
        RECT 31.045 95.665 31.335 96.390 ;
        RECT 31.505 95.665 36.850 96.435 ;
        RECT 37.025 95.665 42.370 96.435 ;
        RECT 42.545 95.665 45.135 96.435 ;
        RECT 45.305 95.665 45.595 96.390 ;
        RECT 45.765 95.665 51.110 96.435 ;
        RECT 51.285 95.665 56.630 96.435 ;
        RECT 56.805 95.665 59.395 96.435 ;
        RECT 59.565 95.665 59.855 96.390 ;
        RECT 60.025 95.665 65.370 96.435 ;
        RECT 65.545 95.665 70.890 96.435 ;
        RECT 71.065 95.665 73.655 96.435 ;
        RECT 73.825 95.665 74.115 96.390 ;
        RECT 74.285 95.665 79.630 96.435 ;
        RECT 79.805 95.665 85.150 96.435 ;
        RECT 85.325 95.665 87.915 96.435 ;
        RECT 88.085 95.665 88.375 96.390 ;
        RECT 88.545 95.665 93.890 96.435 ;
        RECT 94.065 95.665 97.575 96.435 ;
        RECT 99.355 96.415 99.875 96.955 ;
        RECT 98.665 95.665 99.875 96.415 ;
        RECT 16.700 95.495 16.845 95.665 ;
        RECT 17.015 95.495 17.305 95.665 ;
        RECT 17.475 95.495 17.765 95.665 ;
        RECT 17.935 95.495 18.225 95.665 ;
        RECT 18.395 95.495 18.685 95.665 ;
        RECT 18.855 95.495 19.145 95.665 ;
        RECT 19.315 95.495 19.605 95.665 ;
        RECT 19.775 95.495 20.065 95.665 ;
        RECT 20.235 95.495 20.525 95.665 ;
        RECT 20.695 95.495 20.985 95.665 ;
        RECT 21.155 95.495 21.445 95.665 ;
        RECT 21.615 95.495 21.905 95.665 ;
        RECT 22.075 95.495 22.365 95.665 ;
        RECT 22.535 95.495 22.825 95.665 ;
        RECT 22.995 95.495 23.285 95.665 ;
        RECT 23.455 95.495 23.745 95.665 ;
        RECT 23.915 95.495 24.205 95.665 ;
        RECT 24.375 95.495 24.665 95.665 ;
        RECT 24.835 95.495 25.125 95.665 ;
        RECT 25.295 95.495 25.585 95.665 ;
        RECT 25.755 95.495 26.045 95.665 ;
        RECT 26.215 95.495 26.505 95.665 ;
        RECT 26.675 95.495 26.965 95.665 ;
        RECT 27.135 95.495 27.425 95.665 ;
        RECT 27.595 95.495 27.885 95.665 ;
        RECT 28.055 95.495 28.345 95.665 ;
        RECT 28.515 95.495 28.805 95.665 ;
        RECT 28.975 95.495 29.265 95.665 ;
        RECT 29.435 95.495 29.725 95.665 ;
        RECT 29.895 95.495 30.185 95.665 ;
        RECT 30.355 95.495 30.645 95.665 ;
        RECT 30.815 95.495 31.105 95.665 ;
        RECT 31.275 95.495 31.565 95.665 ;
        RECT 31.735 95.495 32.025 95.665 ;
        RECT 32.195 95.495 32.485 95.665 ;
        RECT 32.655 95.495 32.945 95.665 ;
        RECT 33.115 95.495 33.405 95.665 ;
        RECT 33.575 95.495 33.865 95.665 ;
        RECT 34.035 95.495 34.325 95.665 ;
        RECT 34.495 95.495 34.785 95.665 ;
        RECT 34.955 95.495 35.245 95.665 ;
        RECT 35.415 95.495 35.705 95.665 ;
        RECT 35.875 95.495 36.165 95.665 ;
        RECT 36.335 95.495 36.625 95.665 ;
        RECT 36.795 95.495 37.085 95.665 ;
        RECT 37.255 95.495 37.545 95.665 ;
        RECT 37.715 95.495 38.005 95.665 ;
        RECT 38.175 95.495 38.465 95.665 ;
        RECT 38.635 95.495 38.925 95.665 ;
        RECT 39.095 95.495 39.385 95.665 ;
        RECT 39.555 95.495 39.845 95.665 ;
        RECT 40.015 95.495 40.305 95.665 ;
        RECT 40.475 95.495 40.765 95.665 ;
        RECT 40.935 95.495 41.225 95.665 ;
        RECT 41.395 95.495 41.685 95.665 ;
        RECT 41.855 95.495 42.145 95.665 ;
        RECT 42.315 95.495 42.605 95.665 ;
        RECT 42.775 95.495 43.065 95.665 ;
        RECT 43.235 95.495 43.525 95.665 ;
        RECT 43.695 95.495 43.985 95.665 ;
        RECT 44.155 95.495 44.445 95.665 ;
        RECT 44.615 95.495 44.905 95.665 ;
        RECT 45.075 95.495 45.365 95.665 ;
        RECT 45.535 95.495 45.825 95.665 ;
        RECT 45.995 95.495 46.285 95.665 ;
        RECT 46.455 95.495 46.745 95.665 ;
        RECT 46.915 95.495 47.205 95.665 ;
        RECT 47.375 95.495 47.665 95.665 ;
        RECT 47.835 95.495 48.125 95.665 ;
        RECT 48.295 95.495 48.585 95.665 ;
        RECT 48.755 95.495 49.045 95.665 ;
        RECT 49.215 95.495 49.505 95.665 ;
        RECT 49.675 95.495 49.965 95.665 ;
        RECT 50.135 95.495 50.425 95.665 ;
        RECT 50.595 95.495 50.885 95.665 ;
        RECT 51.055 95.495 51.345 95.665 ;
        RECT 51.515 95.495 51.805 95.665 ;
        RECT 51.975 95.495 52.265 95.665 ;
        RECT 52.435 95.495 52.725 95.665 ;
        RECT 52.895 95.495 53.185 95.665 ;
        RECT 53.355 95.495 53.645 95.665 ;
        RECT 53.815 95.495 54.105 95.665 ;
        RECT 54.275 95.495 54.565 95.665 ;
        RECT 54.735 95.495 55.025 95.665 ;
        RECT 55.195 95.495 55.485 95.665 ;
        RECT 55.655 95.495 55.945 95.665 ;
        RECT 56.115 95.495 56.405 95.665 ;
        RECT 56.575 95.495 56.865 95.665 ;
        RECT 57.035 95.495 57.325 95.665 ;
        RECT 57.495 95.495 57.785 95.665 ;
        RECT 57.955 95.495 58.245 95.665 ;
        RECT 58.415 95.495 58.705 95.665 ;
        RECT 58.875 95.495 59.165 95.665 ;
        RECT 59.335 95.495 59.625 95.665 ;
        RECT 59.795 95.495 60.085 95.665 ;
        RECT 60.255 95.495 60.545 95.665 ;
        RECT 60.715 95.495 61.005 95.665 ;
        RECT 61.175 95.495 61.465 95.665 ;
        RECT 61.635 95.495 61.925 95.665 ;
        RECT 62.095 95.495 62.385 95.665 ;
        RECT 62.555 95.495 62.845 95.665 ;
        RECT 63.015 95.495 63.305 95.665 ;
        RECT 63.475 95.495 63.765 95.665 ;
        RECT 63.935 95.495 64.225 95.665 ;
        RECT 64.395 95.495 64.685 95.665 ;
        RECT 64.855 95.495 65.145 95.665 ;
        RECT 65.315 95.495 65.605 95.665 ;
        RECT 65.775 95.495 66.065 95.665 ;
        RECT 66.235 95.495 66.525 95.665 ;
        RECT 66.695 95.495 66.985 95.665 ;
        RECT 67.155 95.495 67.445 95.665 ;
        RECT 67.615 95.495 67.905 95.665 ;
        RECT 68.075 95.495 68.365 95.665 ;
        RECT 68.535 95.495 68.825 95.665 ;
        RECT 68.995 95.495 69.285 95.665 ;
        RECT 69.455 95.495 69.745 95.665 ;
        RECT 69.915 95.495 70.205 95.665 ;
        RECT 70.375 95.495 70.665 95.665 ;
        RECT 70.835 95.495 71.125 95.665 ;
        RECT 71.295 95.495 71.585 95.665 ;
        RECT 71.755 95.495 72.045 95.665 ;
        RECT 72.215 95.495 72.505 95.665 ;
        RECT 72.675 95.495 72.965 95.665 ;
        RECT 73.135 95.495 73.425 95.665 ;
        RECT 73.595 95.495 73.885 95.665 ;
        RECT 74.055 95.495 74.345 95.665 ;
        RECT 74.515 95.495 74.805 95.665 ;
        RECT 74.975 95.495 75.265 95.665 ;
        RECT 75.435 95.495 75.725 95.665 ;
        RECT 75.895 95.495 76.185 95.665 ;
        RECT 76.355 95.495 76.645 95.665 ;
        RECT 76.815 95.495 77.105 95.665 ;
        RECT 77.275 95.495 77.565 95.665 ;
        RECT 77.735 95.495 78.025 95.665 ;
        RECT 78.195 95.495 78.485 95.665 ;
        RECT 78.655 95.495 78.945 95.665 ;
        RECT 79.115 95.495 79.405 95.665 ;
        RECT 79.575 95.495 79.865 95.665 ;
        RECT 80.035 95.495 80.325 95.665 ;
        RECT 80.495 95.495 80.785 95.665 ;
        RECT 80.955 95.495 81.245 95.665 ;
        RECT 81.415 95.495 81.705 95.665 ;
        RECT 81.875 95.495 82.165 95.665 ;
        RECT 82.335 95.495 82.625 95.665 ;
        RECT 82.795 95.495 83.085 95.665 ;
        RECT 83.255 95.495 83.545 95.665 ;
        RECT 83.715 95.495 84.005 95.665 ;
        RECT 84.175 95.495 84.465 95.665 ;
        RECT 84.635 95.495 84.925 95.665 ;
        RECT 85.095 95.495 85.385 95.665 ;
        RECT 85.555 95.495 85.845 95.665 ;
        RECT 86.015 95.495 86.305 95.665 ;
        RECT 86.475 95.495 86.765 95.665 ;
        RECT 86.935 95.495 87.225 95.665 ;
        RECT 87.395 95.495 87.685 95.665 ;
        RECT 87.855 95.495 88.145 95.665 ;
        RECT 88.315 95.495 88.605 95.665 ;
        RECT 88.775 95.495 89.065 95.665 ;
        RECT 89.235 95.495 89.525 95.665 ;
        RECT 89.695 95.495 89.985 95.665 ;
        RECT 90.155 95.495 90.445 95.665 ;
        RECT 90.615 95.495 90.905 95.665 ;
        RECT 91.075 95.495 91.365 95.665 ;
        RECT 91.535 95.495 91.825 95.665 ;
        RECT 91.995 95.495 92.285 95.665 ;
        RECT 92.455 95.495 92.745 95.665 ;
        RECT 92.915 95.495 93.205 95.665 ;
        RECT 93.375 95.495 93.665 95.665 ;
        RECT 93.835 95.495 94.125 95.665 ;
        RECT 94.295 95.495 94.585 95.665 ;
        RECT 94.755 95.495 95.045 95.665 ;
        RECT 95.215 95.495 95.505 95.665 ;
        RECT 95.675 95.495 95.965 95.665 ;
        RECT 96.135 95.495 96.425 95.665 ;
        RECT 96.595 95.495 96.885 95.665 ;
        RECT 97.055 95.495 97.345 95.665 ;
        RECT 97.515 95.495 97.805 95.665 ;
        RECT 97.975 95.495 98.265 95.665 ;
        RECT 98.435 95.495 98.725 95.665 ;
        RECT 98.895 95.495 99.185 95.665 ;
        RECT 99.355 95.495 99.645 95.665 ;
        RECT 99.815 95.495 99.960 95.665 ;
        RECT 16.785 94.745 17.995 95.495 ;
        RECT 18.165 94.745 19.375 95.495 ;
        RECT 16.785 94.205 17.305 94.745 ;
        RECT 17.475 94.035 17.995 94.575 ;
        RECT 18.165 94.205 18.685 94.745 ;
        RECT 18.855 94.035 19.375 94.575 ;
        RECT 16.785 92.945 17.995 94.035 ;
        RECT 18.165 92.945 19.375 94.035 ;
      LAYER li1 ;
        RECT 19.545 93.840 20.065 95.325 ;
      LAYER li1 ;
        RECT 20.235 94.835 20.575 95.495 ;
        RECT 20.925 94.725 26.270 95.495 ;
        RECT 26.445 94.725 29.955 95.495 ;
        RECT 31.045 94.770 31.335 95.495 ;
        RECT 20.925 94.205 23.505 94.725 ;
        RECT 23.675 94.035 26.270 94.555 ;
        RECT 26.445 94.205 28.095 94.725 ;
        RECT 28.265 94.035 29.955 94.555 ;
        RECT 19.735 92.945 20.065 93.670 ;
        RECT 20.925 92.945 26.270 94.035 ;
        RECT 26.445 92.945 29.955 94.035 ;
        RECT 31.045 92.945 31.335 94.110 ;
      LAYER li1 ;
        RECT 31.505 93.840 32.025 95.325 ;
      LAYER li1 ;
        RECT 32.195 94.835 32.535 95.495 ;
        RECT 32.885 94.725 38.230 95.495 ;
        RECT 38.405 94.725 43.750 95.495 ;
        RECT 43.925 94.725 49.270 95.495 ;
        RECT 49.445 94.725 54.790 95.495 ;
        RECT 54.965 94.725 58.475 95.495 ;
        RECT 59.105 94.770 59.395 95.495 ;
        RECT 32.885 94.205 35.465 94.725 ;
        RECT 35.635 94.035 38.230 94.555 ;
        RECT 38.405 94.205 40.985 94.725 ;
        RECT 41.155 94.035 43.750 94.555 ;
        RECT 43.925 94.205 46.505 94.725 ;
        RECT 46.675 94.035 49.270 94.555 ;
        RECT 49.445 94.205 52.025 94.725 ;
        RECT 52.195 94.035 54.790 94.555 ;
        RECT 54.965 94.205 56.615 94.725 ;
        RECT 56.785 94.035 58.475 94.555 ;
        RECT 31.695 92.945 32.025 93.670 ;
        RECT 32.885 92.945 38.230 94.035 ;
        RECT 38.405 92.945 43.750 94.035 ;
        RECT 43.925 92.945 49.270 94.035 ;
        RECT 49.445 92.945 54.790 94.035 ;
        RECT 54.965 92.945 58.475 94.035 ;
        RECT 59.105 92.945 59.395 94.110 ;
      LAYER li1 ;
        RECT 59.565 93.840 60.085 95.325 ;
      LAYER li1 ;
        RECT 60.255 94.835 60.595 95.495 ;
        RECT 60.945 94.725 66.290 95.495 ;
        RECT 66.465 94.725 71.810 95.495 ;
        RECT 71.985 94.725 77.330 95.495 ;
        RECT 77.505 94.725 82.850 95.495 ;
        RECT 83.025 94.725 86.535 95.495 ;
        RECT 87.165 94.770 87.455 95.495 ;
        RECT 60.945 94.205 63.525 94.725 ;
        RECT 63.695 94.035 66.290 94.555 ;
        RECT 66.465 94.205 69.045 94.725 ;
        RECT 69.215 94.035 71.810 94.555 ;
        RECT 71.985 94.205 74.565 94.725 ;
        RECT 74.735 94.035 77.330 94.555 ;
        RECT 77.505 94.205 80.085 94.725 ;
        RECT 80.255 94.035 82.850 94.555 ;
        RECT 83.025 94.205 84.675 94.725 ;
        RECT 84.845 94.035 86.535 94.555 ;
        RECT 59.755 92.945 60.085 93.670 ;
        RECT 60.945 92.945 66.290 94.035 ;
        RECT 66.465 92.945 71.810 94.035 ;
        RECT 71.985 92.945 77.330 94.035 ;
        RECT 77.505 92.945 82.850 94.035 ;
        RECT 83.025 92.945 86.535 94.035 ;
        RECT 87.165 92.945 87.455 94.110 ;
      LAYER li1 ;
        RECT 87.625 93.840 88.145 95.325 ;
      LAYER li1 ;
        RECT 88.315 94.835 88.655 95.495 ;
        RECT 89.005 94.725 92.515 95.495 ;
        RECT 89.005 94.205 90.655 94.725 ;
        RECT 90.825 94.035 92.515 94.555 ;
        RECT 87.815 92.945 88.145 93.670 ;
        RECT 89.005 92.945 92.515 94.035 ;
      LAYER li1 ;
        RECT 93.605 93.840 94.125 95.325 ;
      LAYER li1 ;
        RECT 94.295 94.835 94.635 95.495 ;
        RECT 94.985 94.725 98.495 95.495 ;
        RECT 98.665 94.745 99.875 95.495 ;
        RECT 94.985 94.205 96.635 94.725 ;
        RECT 96.805 94.035 98.495 94.555 ;
        RECT 93.795 92.945 94.125 93.670 ;
        RECT 94.985 92.945 98.495 94.035 ;
        RECT 98.665 94.035 99.185 94.575 ;
        RECT 99.355 94.205 99.875 94.745 ;
        RECT 98.665 92.945 99.875 94.035 ;
        RECT 16.700 92.775 16.845 92.945 ;
        RECT 17.015 92.775 17.305 92.945 ;
        RECT 17.475 92.775 17.765 92.945 ;
        RECT 17.935 92.775 18.225 92.945 ;
        RECT 18.395 92.775 18.685 92.945 ;
        RECT 18.855 92.775 19.145 92.945 ;
        RECT 19.315 92.775 19.605 92.945 ;
        RECT 19.775 92.775 20.065 92.945 ;
        RECT 20.235 92.775 20.525 92.945 ;
        RECT 20.695 92.775 20.985 92.945 ;
        RECT 21.155 92.775 21.445 92.945 ;
        RECT 21.615 92.775 21.905 92.945 ;
        RECT 22.075 92.775 22.365 92.945 ;
        RECT 22.535 92.775 22.825 92.945 ;
        RECT 22.995 92.775 23.285 92.945 ;
        RECT 23.455 92.775 23.745 92.945 ;
        RECT 23.915 92.775 24.205 92.945 ;
        RECT 24.375 92.775 24.665 92.945 ;
        RECT 24.835 92.775 25.125 92.945 ;
        RECT 25.295 92.775 25.585 92.945 ;
        RECT 25.755 92.775 26.045 92.945 ;
        RECT 26.215 92.775 26.505 92.945 ;
        RECT 26.675 92.775 26.965 92.945 ;
        RECT 27.135 92.775 27.425 92.945 ;
        RECT 27.595 92.775 27.885 92.945 ;
        RECT 28.055 92.775 28.345 92.945 ;
        RECT 28.515 92.775 28.805 92.945 ;
        RECT 28.975 92.775 29.265 92.945 ;
        RECT 29.435 92.775 29.725 92.945 ;
        RECT 29.895 92.775 30.185 92.945 ;
        RECT 30.355 92.775 30.645 92.945 ;
        RECT 30.815 92.775 31.105 92.945 ;
        RECT 31.275 92.775 31.565 92.945 ;
        RECT 31.735 92.775 32.025 92.945 ;
        RECT 32.195 92.775 32.485 92.945 ;
        RECT 32.655 92.775 32.945 92.945 ;
        RECT 33.115 92.775 33.405 92.945 ;
        RECT 33.575 92.775 33.865 92.945 ;
        RECT 34.035 92.775 34.325 92.945 ;
        RECT 34.495 92.775 34.785 92.945 ;
        RECT 34.955 92.775 35.245 92.945 ;
        RECT 35.415 92.775 35.705 92.945 ;
        RECT 35.875 92.775 36.165 92.945 ;
        RECT 36.335 92.775 36.625 92.945 ;
        RECT 36.795 92.775 37.085 92.945 ;
        RECT 37.255 92.775 37.545 92.945 ;
        RECT 37.715 92.775 38.005 92.945 ;
        RECT 38.175 92.775 38.465 92.945 ;
        RECT 38.635 92.775 38.925 92.945 ;
        RECT 39.095 92.775 39.385 92.945 ;
        RECT 39.555 92.775 39.845 92.945 ;
        RECT 40.015 92.775 40.305 92.945 ;
        RECT 40.475 92.775 40.765 92.945 ;
        RECT 40.935 92.775 41.225 92.945 ;
        RECT 41.395 92.775 41.685 92.945 ;
        RECT 41.855 92.775 42.145 92.945 ;
        RECT 42.315 92.775 42.605 92.945 ;
        RECT 42.775 92.775 43.065 92.945 ;
        RECT 43.235 92.775 43.525 92.945 ;
        RECT 43.695 92.775 43.985 92.945 ;
        RECT 44.155 92.775 44.445 92.945 ;
        RECT 44.615 92.775 44.905 92.945 ;
        RECT 45.075 92.775 45.365 92.945 ;
        RECT 45.535 92.775 45.825 92.945 ;
        RECT 45.995 92.775 46.285 92.945 ;
        RECT 46.455 92.775 46.745 92.945 ;
        RECT 46.915 92.775 47.205 92.945 ;
        RECT 47.375 92.775 47.665 92.945 ;
        RECT 47.835 92.775 48.125 92.945 ;
        RECT 48.295 92.775 48.585 92.945 ;
        RECT 48.755 92.775 49.045 92.945 ;
        RECT 49.215 92.775 49.505 92.945 ;
        RECT 49.675 92.775 49.965 92.945 ;
        RECT 50.135 92.775 50.425 92.945 ;
        RECT 50.595 92.775 50.885 92.945 ;
        RECT 51.055 92.775 51.345 92.945 ;
        RECT 51.515 92.775 51.805 92.945 ;
        RECT 51.975 92.775 52.265 92.945 ;
        RECT 52.435 92.775 52.725 92.945 ;
        RECT 52.895 92.775 53.185 92.945 ;
        RECT 53.355 92.775 53.645 92.945 ;
        RECT 53.815 92.775 54.105 92.945 ;
        RECT 54.275 92.775 54.565 92.945 ;
        RECT 54.735 92.775 55.025 92.945 ;
        RECT 55.195 92.775 55.485 92.945 ;
        RECT 55.655 92.775 55.945 92.945 ;
        RECT 56.115 92.775 56.405 92.945 ;
        RECT 56.575 92.775 56.865 92.945 ;
        RECT 57.035 92.775 57.325 92.945 ;
        RECT 57.495 92.775 57.785 92.945 ;
        RECT 57.955 92.775 58.245 92.945 ;
        RECT 58.415 92.775 58.705 92.945 ;
        RECT 58.875 92.775 59.165 92.945 ;
        RECT 59.335 92.775 59.625 92.945 ;
        RECT 59.795 92.775 60.085 92.945 ;
        RECT 60.255 92.775 60.545 92.945 ;
        RECT 60.715 92.775 61.005 92.945 ;
        RECT 61.175 92.775 61.465 92.945 ;
        RECT 61.635 92.775 61.925 92.945 ;
        RECT 62.095 92.775 62.385 92.945 ;
        RECT 62.555 92.775 62.845 92.945 ;
        RECT 63.015 92.775 63.305 92.945 ;
        RECT 63.475 92.775 63.765 92.945 ;
        RECT 63.935 92.775 64.225 92.945 ;
        RECT 64.395 92.775 64.685 92.945 ;
        RECT 64.855 92.775 65.145 92.945 ;
        RECT 65.315 92.775 65.605 92.945 ;
        RECT 65.775 92.775 66.065 92.945 ;
        RECT 66.235 92.775 66.525 92.945 ;
        RECT 66.695 92.775 66.985 92.945 ;
        RECT 67.155 92.775 67.445 92.945 ;
        RECT 67.615 92.775 67.905 92.945 ;
        RECT 68.075 92.775 68.365 92.945 ;
        RECT 68.535 92.775 68.825 92.945 ;
        RECT 68.995 92.775 69.285 92.945 ;
        RECT 69.455 92.775 69.745 92.945 ;
        RECT 69.915 92.775 70.205 92.945 ;
        RECT 70.375 92.775 70.665 92.945 ;
        RECT 70.835 92.775 71.125 92.945 ;
        RECT 71.295 92.775 71.585 92.945 ;
        RECT 71.755 92.775 72.045 92.945 ;
        RECT 72.215 92.775 72.505 92.945 ;
        RECT 72.675 92.775 72.965 92.945 ;
        RECT 73.135 92.775 73.425 92.945 ;
        RECT 73.595 92.775 73.885 92.945 ;
        RECT 74.055 92.775 74.345 92.945 ;
        RECT 74.515 92.775 74.805 92.945 ;
        RECT 74.975 92.775 75.265 92.945 ;
        RECT 75.435 92.775 75.725 92.945 ;
        RECT 75.895 92.775 76.185 92.945 ;
        RECT 76.355 92.775 76.645 92.945 ;
        RECT 76.815 92.775 77.105 92.945 ;
        RECT 77.275 92.775 77.565 92.945 ;
        RECT 77.735 92.775 78.025 92.945 ;
        RECT 78.195 92.775 78.485 92.945 ;
        RECT 78.655 92.775 78.945 92.945 ;
        RECT 79.115 92.775 79.405 92.945 ;
        RECT 79.575 92.775 79.865 92.945 ;
        RECT 80.035 92.775 80.325 92.945 ;
        RECT 80.495 92.775 80.785 92.945 ;
        RECT 80.955 92.775 81.245 92.945 ;
        RECT 81.415 92.775 81.705 92.945 ;
        RECT 81.875 92.775 82.165 92.945 ;
        RECT 82.335 92.775 82.625 92.945 ;
        RECT 82.795 92.775 83.085 92.945 ;
        RECT 83.255 92.775 83.545 92.945 ;
        RECT 83.715 92.775 84.005 92.945 ;
        RECT 84.175 92.775 84.465 92.945 ;
        RECT 84.635 92.775 84.925 92.945 ;
        RECT 85.095 92.775 85.385 92.945 ;
        RECT 85.555 92.775 85.845 92.945 ;
        RECT 86.015 92.775 86.305 92.945 ;
        RECT 86.475 92.775 86.765 92.945 ;
        RECT 86.935 92.775 87.225 92.945 ;
        RECT 87.395 92.775 87.685 92.945 ;
        RECT 87.855 92.775 88.145 92.945 ;
        RECT 88.315 92.775 88.605 92.945 ;
        RECT 88.775 92.775 89.065 92.945 ;
        RECT 89.235 92.775 89.525 92.945 ;
        RECT 89.695 92.775 89.985 92.945 ;
        RECT 90.155 92.775 90.445 92.945 ;
        RECT 90.615 92.775 90.905 92.945 ;
        RECT 91.075 92.775 91.365 92.945 ;
        RECT 91.535 92.775 91.825 92.945 ;
        RECT 91.995 92.775 92.285 92.945 ;
        RECT 92.455 92.775 92.745 92.945 ;
        RECT 92.915 92.775 93.205 92.945 ;
        RECT 93.375 92.775 93.665 92.945 ;
        RECT 93.835 92.775 94.125 92.945 ;
        RECT 94.295 92.775 94.585 92.945 ;
        RECT 94.755 92.775 95.045 92.945 ;
        RECT 95.215 92.775 95.505 92.945 ;
        RECT 95.675 92.775 95.965 92.945 ;
        RECT 96.135 92.775 96.425 92.945 ;
        RECT 96.595 92.775 96.885 92.945 ;
        RECT 97.055 92.775 97.345 92.945 ;
        RECT 97.515 92.775 97.805 92.945 ;
        RECT 97.975 92.775 98.265 92.945 ;
        RECT 98.435 92.775 98.725 92.945 ;
        RECT 98.895 92.775 99.185 92.945 ;
        RECT 99.355 92.775 99.645 92.945 ;
        RECT 99.815 92.775 99.960 92.945 ;
        RECT 16.785 91.685 17.995 92.775 ;
        RECT 18.165 91.685 23.510 92.775 ;
        RECT 23.685 91.685 29.030 92.775 ;
        RECT 29.205 91.685 34.550 92.775 ;
        RECT 34.725 91.685 40.070 92.775 ;
        RECT 40.245 91.685 43.755 92.775 ;
        RECT 16.785 90.975 17.305 91.515 ;
        RECT 17.475 91.145 17.995 91.685 ;
        RECT 18.165 90.995 20.745 91.515 ;
        RECT 20.915 91.165 23.510 91.685 ;
        RECT 23.685 90.995 26.265 91.515 ;
        RECT 26.435 91.165 29.030 91.685 ;
        RECT 29.205 90.995 31.785 91.515 ;
        RECT 31.955 91.165 34.550 91.685 ;
        RECT 34.725 90.995 37.305 91.515 ;
        RECT 37.475 91.165 40.070 91.685 ;
        RECT 40.245 90.995 41.895 91.515 ;
        RECT 42.065 91.165 43.755 91.685 ;
        RECT 44.845 91.610 45.135 92.775 ;
        RECT 45.305 91.685 50.650 92.775 ;
        RECT 50.825 91.685 56.170 92.775 ;
        RECT 56.345 91.685 61.690 92.775 ;
        RECT 61.865 91.685 63.535 92.775 ;
        RECT 64.175 92.020 64.505 92.775 ;
        RECT 64.685 91.890 64.865 92.605 ;
        RECT 65.070 92.075 65.400 92.775 ;
      LAYER li1 ;
        RECT 65.610 91.900 65.800 92.605 ;
      LAYER li1 ;
        RECT 65.970 92.075 66.300 92.775 ;
      LAYER li1 ;
        RECT 66.470 91.905 66.660 92.605 ;
      LAYER li1 ;
        RECT 66.830 92.075 67.160 92.775 ;
      LAYER li1 ;
        RECT 66.470 91.900 67.215 91.905 ;
      LAYER li1 ;
        RECT 45.305 90.995 47.885 91.515 ;
        RECT 48.055 91.165 50.650 91.685 ;
        RECT 50.825 90.995 53.405 91.515 ;
        RECT 53.575 91.165 56.170 91.685 ;
        RECT 56.345 90.995 58.925 91.515 ;
        RECT 59.095 91.165 61.690 91.685 ;
        RECT 61.865 90.995 62.615 91.515 ;
        RECT 62.785 91.165 63.535 91.685 ;
      LAYER li1 ;
        RECT 64.205 91.135 64.515 91.755 ;
      LAYER li1 ;
        RECT 64.685 91.720 65.440 91.890 ;
        RECT 65.230 91.495 65.440 91.720 ;
      LAYER li1 ;
        RECT 65.610 91.675 67.215 91.900 ;
      LAYER li1 ;
        RECT 67.385 91.685 72.730 92.775 ;
        RECT 65.230 91.160 66.765 91.495 ;
        RECT 16.785 90.225 17.995 90.975 ;
        RECT 18.165 90.225 23.510 90.995 ;
        RECT 23.685 90.225 29.030 90.995 ;
        RECT 29.205 90.225 34.550 90.995 ;
        RECT 34.725 90.225 40.070 90.995 ;
        RECT 40.245 90.225 43.755 90.995 ;
        RECT 44.845 90.225 45.135 90.950 ;
        RECT 45.305 90.225 50.650 90.995 ;
        RECT 50.825 90.225 56.170 90.995 ;
        RECT 56.345 90.225 61.690 90.995 ;
        RECT 61.865 90.225 63.535 90.995 ;
        RECT 65.230 90.945 65.440 91.160 ;
      LAYER li1 ;
        RECT 66.935 90.985 67.215 91.675 ;
      LAYER li1 ;
        RECT 64.175 90.755 65.440 90.945 ;
      LAYER li1 ;
        RECT 65.610 90.755 67.215 90.985 ;
      LAYER li1 ;
        RECT 67.385 90.995 69.965 91.515 ;
        RECT 70.135 91.165 72.730 91.685 ;
        RECT 72.905 91.610 73.195 92.775 ;
        RECT 73.365 91.685 78.710 92.775 ;
        RECT 78.885 91.685 84.230 92.775 ;
        RECT 84.405 91.685 89.750 92.775 ;
        RECT 89.925 91.685 93.435 92.775 ;
        RECT 93.795 92.050 94.125 92.775 ;
        RECT 73.365 90.995 75.945 91.515 ;
        RECT 76.115 91.165 78.710 91.685 ;
        RECT 78.885 90.995 81.465 91.515 ;
        RECT 81.635 91.165 84.230 91.685 ;
        RECT 84.405 90.995 86.985 91.515 ;
        RECT 87.155 91.165 89.750 91.685 ;
        RECT 89.925 90.995 91.575 91.515 ;
        RECT 91.745 91.165 93.435 91.685 ;
        RECT 64.175 90.395 64.505 90.755 ;
      LAYER li1 ;
        RECT 65.610 90.655 65.800 90.755 ;
      LAYER li1 ;
        RECT 65.035 90.225 65.365 90.585 ;
        RECT 65.970 90.225 66.300 90.585 ;
      LAYER li1 ;
        RECT 66.470 90.395 66.660 90.755 ;
      LAYER li1 ;
        RECT 66.830 90.225 67.160 90.585 ;
        RECT 67.385 90.225 72.730 90.995 ;
        RECT 72.905 90.225 73.195 90.950 ;
        RECT 73.365 90.225 78.710 90.995 ;
        RECT 78.885 90.225 84.230 90.995 ;
        RECT 84.405 90.225 89.750 90.995 ;
        RECT 89.925 90.225 93.435 90.995 ;
      LAYER li1 ;
        RECT 93.605 90.395 94.125 91.880 ;
      LAYER li1 ;
        RECT 94.985 91.685 98.495 92.775 ;
        RECT 94.985 90.995 96.635 91.515 ;
        RECT 96.805 91.165 98.495 91.685 ;
        RECT 98.665 91.685 99.875 92.775 ;
        RECT 98.665 91.145 99.185 91.685 ;
        RECT 94.295 90.225 94.635 90.885 ;
        RECT 94.985 90.225 98.495 90.995 ;
        RECT 99.355 90.975 99.875 91.515 ;
        RECT 98.665 90.225 99.875 90.975 ;
        RECT 16.700 90.055 16.845 90.225 ;
        RECT 17.015 90.055 17.305 90.225 ;
        RECT 17.475 90.055 17.765 90.225 ;
        RECT 17.935 90.055 18.225 90.225 ;
        RECT 18.395 90.055 18.685 90.225 ;
        RECT 18.855 90.055 19.145 90.225 ;
        RECT 19.315 90.055 19.605 90.225 ;
        RECT 19.775 90.055 20.065 90.225 ;
        RECT 20.235 90.055 20.525 90.225 ;
        RECT 20.695 90.055 20.985 90.225 ;
        RECT 21.155 90.055 21.445 90.225 ;
        RECT 21.615 90.055 21.905 90.225 ;
        RECT 22.075 90.055 22.365 90.225 ;
        RECT 22.535 90.055 22.825 90.225 ;
        RECT 22.995 90.055 23.285 90.225 ;
        RECT 23.455 90.055 23.745 90.225 ;
        RECT 23.915 90.055 24.205 90.225 ;
        RECT 24.375 90.055 24.665 90.225 ;
        RECT 24.835 90.055 25.125 90.225 ;
        RECT 25.295 90.055 25.585 90.225 ;
        RECT 25.755 90.055 26.045 90.225 ;
        RECT 26.215 90.055 26.505 90.225 ;
        RECT 26.675 90.055 26.965 90.225 ;
        RECT 27.135 90.055 27.425 90.225 ;
        RECT 27.595 90.055 27.885 90.225 ;
        RECT 28.055 90.055 28.345 90.225 ;
        RECT 28.515 90.055 28.805 90.225 ;
        RECT 28.975 90.055 29.265 90.225 ;
        RECT 29.435 90.055 29.725 90.225 ;
        RECT 29.895 90.055 30.185 90.225 ;
        RECT 30.355 90.055 30.645 90.225 ;
        RECT 30.815 90.055 31.105 90.225 ;
        RECT 31.275 90.055 31.565 90.225 ;
        RECT 31.735 90.055 32.025 90.225 ;
        RECT 32.195 90.055 32.485 90.225 ;
        RECT 32.655 90.055 32.945 90.225 ;
        RECT 33.115 90.055 33.405 90.225 ;
        RECT 33.575 90.055 33.865 90.225 ;
        RECT 34.035 90.055 34.325 90.225 ;
        RECT 34.495 90.055 34.785 90.225 ;
        RECT 34.955 90.055 35.245 90.225 ;
        RECT 35.415 90.055 35.705 90.225 ;
        RECT 35.875 90.055 36.165 90.225 ;
        RECT 36.335 90.055 36.625 90.225 ;
        RECT 36.795 90.055 37.085 90.225 ;
        RECT 37.255 90.055 37.545 90.225 ;
        RECT 37.715 90.055 38.005 90.225 ;
        RECT 38.175 90.055 38.465 90.225 ;
        RECT 38.635 90.055 38.925 90.225 ;
        RECT 39.095 90.055 39.385 90.225 ;
        RECT 39.555 90.055 39.845 90.225 ;
        RECT 40.015 90.055 40.305 90.225 ;
        RECT 40.475 90.055 40.765 90.225 ;
        RECT 40.935 90.055 41.225 90.225 ;
        RECT 41.395 90.055 41.685 90.225 ;
        RECT 41.855 90.055 42.145 90.225 ;
        RECT 42.315 90.055 42.605 90.225 ;
        RECT 42.775 90.055 43.065 90.225 ;
        RECT 43.235 90.055 43.525 90.225 ;
        RECT 43.695 90.055 43.985 90.225 ;
        RECT 44.155 90.055 44.445 90.225 ;
        RECT 44.615 90.055 44.905 90.225 ;
        RECT 45.075 90.055 45.365 90.225 ;
        RECT 45.535 90.055 45.825 90.225 ;
        RECT 45.995 90.055 46.285 90.225 ;
        RECT 46.455 90.055 46.745 90.225 ;
        RECT 46.915 90.055 47.205 90.225 ;
        RECT 47.375 90.055 47.665 90.225 ;
        RECT 47.835 90.055 48.125 90.225 ;
        RECT 48.295 90.055 48.585 90.225 ;
        RECT 48.755 90.055 49.045 90.225 ;
        RECT 49.215 90.055 49.505 90.225 ;
        RECT 49.675 90.055 49.965 90.225 ;
        RECT 50.135 90.055 50.425 90.225 ;
        RECT 50.595 90.055 50.885 90.225 ;
        RECT 51.055 90.055 51.345 90.225 ;
        RECT 51.515 90.055 51.805 90.225 ;
        RECT 51.975 90.055 52.265 90.225 ;
        RECT 52.435 90.055 52.725 90.225 ;
        RECT 52.895 90.055 53.185 90.225 ;
        RECT 53.355 90.055 53.645 90.225 ;
        RECT 53.815 90.055 54.105 90.225 ;
        RECT 54.275 90.055 54.565 90.225 ;
        RECT 54.735 90.055 55.025 90.225 ;
        RECT 55.195 90.055 55.485 90.225 ;
        RECT 55.655 90.055 55.945 90.225 ;
        RECT 56.115 90.055 56.405 90.225 ;
        RECT 56.575 90.055 56.865 90.225 ;
        RECT 57.035 90.055 57.325 90.225 ;
        RECT 57.495 90.055 57.785 90.225 ;
        RECT 57.955 90.055 58.245 90.225 ;
        RECT 58.415 90.055 58.705 90.225 ;
        RECT 58.875 90.055 59.165 90.225 ;
        RECT 59.335 90.055 59.625 90.225 ;
        RECT 59.795 90.055 60.085 90.225 ;
        RECT 60.255 90.055 60.545 90.225 ;
        RECT 60.715 90.055 61.005 90.225 ;
        RECT 61.175 90.055 61.465 90.225 ;
        RECT 61.635 90.055 61.925 90.225 ;
        RECT 62.095 90.055 62.385 90.225 ;
        RECT 62.555 90.055 62.845 90.225 ;
        RECT 63.015 90.055 63.305 90.225 ;
        RECT 63.475 90.055 63.765 90.225 ;
        RECT 63.935 90.055 64.225 90.225 ;
        RECT 64.395 90.055 64.685 90.225 ;
        RECT 64.855 90.055 65.145 90.225 ;
        RECT 65.315 90.055 65.605 90.225 ;
        RECT 65.775 90.055 66.065 90.225 ;
        RECT 66.235 90.055 66.525 90.225 ;
        RECT 66.695 90.055 66.985 90.225 ;
        RECT 67.155 90.055 67.445 90.225 ;
        RECT 67.615 90.055 67.905 90.225 ;
        RECT 68.075 90.055 68.365 90.225 ;
        RECT 68.535 90.055 68.825 90.225 ;
        RECT 68.995 90.055 69.285 90.225 ;
        RECT 69.455 90.055 69.745 90.225 ;
        RECT 69.915 90.055 70.205 90.225 ;
        RECT 70.375 90.055 70.665 90.225 ;
        RECT 70.835 90.055 71.125 90.225 ;
        RECT 71.295 90.055 71.585 90.225 ;
        RECT 71.755 90.055 72.045 90.225 ;
        RECT 72.215 90.055 72.505 90.225 ;
        RECT 72.675 90.055 72.965 90.225 ;
        RECT 73.135 90.055 73.425 90.225 ;
        RECT 73.595 90.055 73.885 90.225 ;
        RECT 74.055 90.055 74.345 90.225 ;
        RECT 74.515 90.055 74.805 90.225 ;
        RECT 74.975 90.055 75.265 90.225 ;
        RECT 75.435 90.055 75.725 90.225 ;
        RECT 75.895 90.055 76.185 90.225 ;
        RECT 76.355 90.055 76.645 90.225 ;
        RECT 76.815 90.055 77.105 90.225 ;
        RECT 77.275 90.055 77.565 90.225 ;
        RECT 77.735 90.055 78.025 90.225 ;
        RECT 78.195 90.055 78.485 90.225 ;
        RECT 78.655 90.055 78.945 90.225 ;
        RECT 79.115 90.055 79.405 90.225 ;
        RECT 79.575 90.055 79.865 90.225 ;
        RECT 80.035 90.055 80.325 90.225 ;
        RECT 80.495 90.055 80.785 90.225 ;
        RECT 80.955 90.055 81.245 90.225 ;
        RECT 81.415 90.055 81.705 90.225 ;
        RECT 81.875 90.055 82.165 90.225 ;
        RECT 82.335 90.055 82.625 90.225 ;
        RECT 82.795 90.055 83.085 90.225 ;
        RECT 83.255 90.055 83.545 90.225 ;
        RECT 83.715 90.055 84.005 90.225 ;
        RECT 84.175 90.055 84.465 90.225 ;
        RECT 84.635 90.055 84.925 90.225 ;
        RECT 85.095 90.055 85.385 90.225 ;
        RECT 85.555 90.055 85.845 90.225 ;
        RECT 86.015 90.055 86.305 90.225 ;
        RECT 86.475 90.055 86.765 90.225 ;
        RECT 86.935 90.055 87.225 90.225 ;
        RECT 87.395 90.055 87.685 90.225 ;
        RECT 87.855 90.055 88.145 90.225 ;
        RECT 88.315 90.055 88.605 90.225 ;
        RECT 88.775 90.055 89.065 90.225 ;
        RECT 89.235 90.055 89.525 90.225 ;
        RECT 89.695 90.055 89.985 90.225 ;
        RECT 90.155 90.055 90.445 90.225 ;
        RECT 90.615 90.055 90.905 90.225 ;
        RECT 91.075 90.055 91.365 90.225 ;
        RECT 91.535 90.055 91.825 90.225 ;
        RECT 91.995 90.055 92.285 90.225 ;
        RECT 92.455 90.055 92.745 90.225 ;
        RECT 92.915 90.055 93.205 90.225 ;
        RECT 93.375 90.055 93.665 90.225 ;
        RECT 93.835 90.055 94.125 90.225 ;
        RECT 94.295 90.055 94.585 90.225 ;
        RECT 94.755 90.055 95.045 90.225 ;
        RECT 95.215 90.055 95.505 90.225 ;
        RECT 95.675 90.055 95.965 90.225 ;
        RECT 96.135 90.055 96.425 90.225 ;
        RECT 96.595 90.055 96.885 90.225 ;
        RECT 97.055 90.055 97.345 90.225 ;
        RECT 97.515 90.055 97.805 90.225 ;
        RECT 97.975 90.055 98.265 90.225 ;
        RECT 98.435 90.055 98.725 90.225 ;
        RECT 98.895 90.055 99.185 90.225 ;
        RECT 99.355 90.055 99.645 90.225 ;
        RECT 99.815 90.055 99.960 90.225 ;
        RECT 16.785 89.305 17.995 90.055 ;
        RECT 16.785 88.765 17.305 89.305 ;
        RECT 18.165 89.285 23.510 90.055 ;
        RECT 23.685 89.285 29.030 90.055 ;
        RECT 29.205 89.285 30.875 90.055 ;
        RECT 31.045 89.330 31.335 90.055 ;
        RECT 31.505 89.285 36.850 90.055 ;
        RECT 37.025 89.285 42.370 90.055 ;
        RECT 42.545 89.285 47.890 90.055 ;
        RECT 48.065 89.285 53.410 90.055 ;
        RECT 53.585 89.285 58.930 90.055 ;
        RECT 59.105 89.330 59.395 90.055 ;
        RECT 59.565 89.285 62.155 90.055 ;
        RECT 62.415 89.505 62.585 89.795 ;
        RECT 62.755 89.675 63.085 90.055 ;
        RECT 62.415 89.335 63.080 89.505 ;
        RECT 17.475 88.595 17.995 89.135 ;
        RECT 18.165 88.765 20.745 89.285 ;
        RECT 20.915 88.595 23.510 89.115 ;
        RECT 23.685 88.765 26.265 89.285 ;
        RECT 26.435 88.595 29.030 89.115 ;
        RECT 29.205 88.765 29.955 89.285 ;
        RECT 30.125 88.595 30.875 89.115 ;
        RECT 31.505 88.765 34.085 89.285 ;
        RECT 16.785 87.505 17.995 88.595 ;
        RECT 18.165 87.505 23.510 88.595 ;
        RECT 23.685 87.505 29.030 88.595 ;
        RECT 29.205 87.505 30.875 88.595 ;
        RECT 31.045 87.505 31.335 88.670 ;
        RECT 34.255 88.595 36.850 89.115 ;
        RECT 37.025 88.765 39.605 89.285 ;
        RECT 39.775 88.595 42.370 89.115 ;
        RECT 42.545 88.765 45.125 89.285 ;
        RECT 45.295 88.595 47.890 89.115 ;
        RECT 48.065 88.765 50.645 89.285 ;
        RECT 50.815 88.595 53.410 89.115 ;
        RECT 53.585 88.765 56.165 89.285 ;
        RECT 56.335 88.595 58.930 89.115 ;
        RECT 59.565 88.765 60.775 89.285 ;
        RECT 31.505 87.505 36.850 88.595 ;
        RECT 37.025 87.505 42.370 88.595 ;
        RECT 42.545 87.505 47.890 88.595 ;
        RECT 48.065 87.505 53.410 88.595 ;
        RECT 53.585 87.505 58.930 88.595 ;
        RECT 59.105 87.505 59.395 88.670 ;
        RECT 60.945 88.595 62.155 89.115 ;
        RECT 59.565 87.505 62.155 88.595 ;
      LAYER li1 ;
        RECT 62.330 88.515 62.680 89.165 ;
      LAYER li1 ;
        RECT 62.850 88.345 63.080 89.335 ;
        RECT 62.415 88.175 63.080 88.345 ;
        RECT 62.415 87.675 62.585 88.175 ;
        RECT 62.755 87.505 63.085 88.005 ;
        RECT 63.255 87.675 63.480 89.795 ;
        RECT 63.695 89.595 63.945 90.055 ;
        RECT 64.130 89.605 64.460 89.775 ;
        RECT 64.640 89.605 65.390 89.775 ;
      LAYER li1 ;
        RECT 63.680 88.475 63.960 89.075 ;
      LAYER li1 ;
        RECT 64.130 88.075 64.300 89.605 ;
        RECT 64.470 89.105 65.050 89.435 ;
        RECT 64.470 88.235 64.710 89.105 ;
        RECT 65.220 88.825 65.390 89.605 ;
        RECT 65.640 89.555 66.010 90.055 ;
        RECT 66.190 89.605 66.650 89.775 ;
        RECT 66.880 89.605 67.550 89.775 ;
        RECT 66.190 89.375 66.360 89.605 ;
        RECT 65.560 89.075 66.360 89.375 ;
        RECT 66.530 89.105 67.080 89.435 ;
        RECT 65.560 89.045 65.730 89.075 ;
        RECT 65.850 88.825 66.020 88.895 ;
        RECT 65.220 88.655 66.020 88.825 ;
        RECT 65.510 88.565 66.020 88.655 ;
        RECT 64.900 88.130 65.340 88.485 ;
        RECT 63.680 87.505 63.945 87.965 ;
        RECT 64.130 87.700 64.365 88.075 ;
        RECT 65.510 87.950 65.680 88.565 ;
        RECT 64.610 87.780 65.680 87.950 ;
        RECT 65.850 87.505 66.020 88.305 ;
        RECT 66.190 88.005 66.360 89.075 ;
        RECT 66.530 88.175 66.720 88.895 ;
        RECT 66.890 88.565 67.080 89.105 ;
        RECT 67.380 89.065 67.550 89.605 ;
        RECT 67.865 89.525 68.035 90.055 ;
        RECT 68.330 89.405 68.690 89.845 ;
        RECT 68.865 89.575 69.035 90.055 ;
        RECT 69.735 89.580 69.905 90.055 ;
        RECT 70.585 89.580 70.755 90.055 ;
        RECT 68.330 89.235 68.830 89.405 ;
        RECT 68.660 89.065 68.830 89.235 ;
        RECT 71.065 89.285 76.410 90.055 ;
        RECT 76.585 89.285 81.930 90.055 ;
        RECT 82.105 89.285 85.615 90.055 ;
        RECT 85.785 89.305 86.995 90.055 ;
        RECT 87.165 89.330 87.455 90.055 ;
        RECT 67.380 88.895 68.470 89.065 ;
        RECT 68.660 88.895 70.480 89.065 ;
        RECT 66.890 88.235 67.210 88.565 ;
        RECT 66.190 87.675 66.440 88.005 ;
        RECT 67.380 87.975 67.550 88.895 ;
        RECT 68.660 88.640 68.830 88.895 ;
        RECT 71.065 88.765 73.645 89.285 ;
        RECT 67.720 88.470 68.830 88.640 ;
        RECT 73.815 88.595 76.410 89.115 ;
        RECT 76.585 88.765 79.165 89.285 ;
        RECT 79.335 88.595 81.930 89.115 ;
        RECT 82.105 88.765 83.755 89.285 ;
        RECT 83.925 88.595 85.615 89.115 ;
        RECT 85.785 88.765 86.305 89.305 ;
        RECT 87.625 89.285 92.970 90.055 ;
        RECT 93.145 89.285 98.490 90.055 ;
        RECT 98.665 89.305 99.875 90.055 ;
        RECT 86.475 88.595 86.995 89.135 ;
        RECT 87.625 88.765 90.205 89.285 ;
        RECT 67.720 88.310 68.580 88.470 ;
        RECT 66.665 87.805 67.550 87.975 ;
        RECT 67.730 87.505 67.945 88.005 ;
        RECT 68.410 87.685 68.580 88.310 ;
        RECT 68.865 87.505 69.045 88.285 ;
        RECT 69.740 87.505 69.910 88.335 ;
        RECT 70.580 87.505 70.750 88.335 ;
        RECT 71.065 87.505 76.410 88.595 ;
        RECT 76.585 87.505 81.930 88.595 ;
        RECT 82.105 87.505 85.615 88.595 ;
        RECT 85.785 87.505 86.995 88.595 ;
        RECT 87.165 87.505 87.455 88.670 ;
        RECT 90.375 88.595 92.970 89.115 ;
        RECT 93.145 88.765 95.725 89.285 ;
        RECT 95.895 88.595 98.490 89.115 ;
        RECT 87.625 87.505 92.970 88.595 ;
        RECT 93.145 87.505 98.490 88.595 ;
        RECT 98.665 88.595 99.185 89.135 ;
        RECT 99.355 88.765 99.875 89.305 ;
        RECT 98.665 87.505 99.875 88.595 ;
        RECT 16.700 87.335 16.845 87.505 ;
        RECT 17.015 87.335 17.305 87.505 ;
        RECT 17.475 87.335 17.765 87.505 ;
        RECT 17.935 87.335 18.225 87.505 ;
        RECT 18.395 87.335 18.685 87.505 ;
        RECT 18.855 87.335 19.145 87.505 ;
        RECT 19.315 87.335 19.605 87.505 ;
        RECT 19.775 87.335 20.065 87.505 ;
        RECT 20.235 87.335 20.525 87.505 ;
        RECT 20.695 87.335 20.985 87.505 ;
        RECT 21.155 87.335 21.445 87.505 ;
        RECT 21.615 87.335 21.905 87.505 ;
        RECT 22.075 87.335 22.365 87.505 ;
        RECT 22.535 87.335 22.825 87.505 ;
        RECT 22.995 87.335 23.285 87.505 ;
        RECT 23.455 87.335 23.745 87.505 ;
        RECT 23.915 87.335 24.205 87.505 ;
        RECT 24.375 87.335 24.665 87.505 ;
        RECT 24.835 87.335 25.125 87.505 ;
        RECT 25.295 87.335 25.585 87.505 ;
        RECT 25.755 87.335 26.045 87.505 ;
        RECT 26.215 87.335 26.505 87.505 ;
        RECT 26.675 87.335 26.965 87.505 ;
        RECT 27.135 87.335 27.425 87.505 ;
        RECT 27.595 87.335 27.885 87.505 ;
        RECT 28.055 87.335 28.345 87.505 ;
        RECT 28.515 87.335 28.805 87.505 ;
        RECT 28.975 87.335 29.265 87.505 ;
        RECT 29.435 87.335 29.725 87.505 ;
        RECT 29.895 87.335 30.185 87.505 ;
        RECT 30.355 87.335 30.645 87.505 ;
        RECT 30.815 87.335 31.105 87.505 ;
        RECT 31.275 87.335 31.565 87.505 ;
        RECT 31.735 87.335 32.025 87.505 ;
        RECT 32.195 87.335 32.485 87.505 ;
        RECT 32.655 87.335 32.945 87.505 ;
        RECT 33.115 87.335 33.405 87.505 ;
        RECT 33.575 87.335 33.865 87.505 ;
        RECT 34.035 87.335 34.325 87.505 ;
        RECT 34.495 87.335 34.785 87.505 ;
        RECT 34.955 87.335 35.245 87.505 ;
        RECT 35.415 87.335 35.705 87.505 ;
        RECT 35.875 87.335 36.165 87.505 ;
        RECT 36.335 87.335 36.625 87.505 ;
        RECT 36.795 87.335 37.085 87.505 ;
        RECT 37.255 87.335 37.545 87.505 ;
        RECT 37.715 87.335 38.005 87.505 ;
        RECT 38.175 87.335 38.465 87.505 ;
        RECT 38.635 87.335 38.925 87.505 ;
        RECT 39.095 87.335 39.385 87.505 ;
        RECT 39.555 87.335 39.845 87.505 ;
        RECT 40.015 87.335 40.305 87.505 ;
        RECT 40.475 87.335 40.765 87.505 ;
        RECT 40.935 87.335 41.225 87.505 ;
        RECT 41.395 87.335 41.685 87.505 ;
        RECT 41.855 87.335 42.145 87.505 ;
        RECT 42.315 87.335 42.605 87.505 ;
        RECT 42.775 87.335 43.065 87.505 ;
        RECT 43.235 87.335 43.525 87.505 ;
        RECT 43.695 87.335 43.985 87.505 ;
        RECT 44.155 87.335 44.445 87.505 ;
        RECT 44.615 87.335 44.905 87.505 ;
        RECT 45.075 87.335 45.365 87.505 ;
        RECT 45.535 87.335 45.825 87.505 ;
        RECT 45.995 87.335 46.285 87.505 ;
        RECT 46.455 87.335 46.745 87.505 ;
        RECT 46.915 87.335 47.205 87.505 ;
        RECT 47.375 87.335 47.665 87.505 ;
        RECT 47.835 87.335 48.125 87.505 ;
        RECT 48.295 87.335 48.585 87.505 ;
        RECT 48.755 87.335 49.045 87.505 ;
        RECT 49.215 87.335 49.505 87.505 ;
        RECT 49.675 87.335 49.965 87.505 ;
        RECT 50.135 87.335 50.425 87.505 ;
        RECT 50.595 87.335 50.885 87.505 ;
        RECT 51.055 87.335 51.345 87.505 ;
        RECT 51.515 87.335 51.805 87.505 ;
        RECT 51.975 87.335 52.265 87.505 ;
        RECT 52.435 87.335 52.725 87.505 ;
        RECT 52.895 87.335 53.185 87.505 ;
        RECT 53.355 87.335 53.645 87.505 ;
        RECT 53.815 87.335 54.105 87.505 ;
        RECT 54.275 87.335 54.565 87.505 ;
        RECT 54.735 87.335 55.025 87.505 ;
        RECT 55.195 87.335 55.485 87.505 ;
        RECT 55.655 87.335 55.945 87.505 ;
        RECT 56.115 87.335 56.405 87.505 ;
        RECT 56.575 87.335 56.865 87.505 ;
        RECT 57.035 87.335 57.325 87.505 ;
        RECT 57.495 87.335 57.785 87.505 ;
        RECT 57.955 87.335 58.245 87.505 ;
        RECT 58.415 87.335 58.705 87.505 ;
        RECT 58.875 87.335 59.165 87.505 ;
        RECT 59.335 87.335 59.625 87.505 ;
        RECT 59.795 87.335 60.085 87.505 ;
        RECT 60.255 87.335 60.545 87.505 ;
        RECT 60.715 87.335 61.005 87.505 ;
        RECT 61.175 87.335 61.465 87.505 ;
        RECT 61.635 87.335 61.925 87.505 ;
        RECT 62.095 87.335 62.385 87.505 ;
        RECT 62.555 87.335 62.845 87.505 ;
        RECT 63.015 87.335 63.305 87.505 ;
        RECT 63.475 87.335 63.765 87.505 ;
        RECT 63.935 87.335 64.225 87.505 ;
        RECT 64.395 87.335 64.685 87.505 ;
        RECT 64.855 87.335 65.145 87.505 ;
        RECT 65.315 87.335 65.605 87.505 ;
        RECT 65.775 87.335 66.065 87.505 ;
        RECT 66.235 87.335 66.525 87.505 ;
        RECT 66.695 87.335 66.985 87.505 ;
        RECT 67.155 87.335 67.445 87.505 ;
        RECT 67.615 87.335 67.905 87.505 ;
        RECT 68.075 87.335 68.365 87.505 ;
        RECT 68.535 87.335 68.825 87.505 ;
        RECT 68.995 87.335 69.285 87.505 ;
        RECT 69.455 87.335 69.745 87.505 ;
        RECT 69.915 87.335 70.205 87.505 ;
        RECT 70.375 87.335 70.665 87.505 ;
        RECT 70.835 87.335 71.125 87.505 ;
        RECT 71.295 87.335 71.585 87.505 ;
        RECT 71.755 87.335 72.045 87.505 ;
        RECT 72.215 87.335 72.505 87.505 ;
        RECT 72.675 87.335 72.965 87.505 ;
        RECT 73.135 87.335 73.425 87.505 ;
        RECT 73.595 87.335 73.885 87.505 ;
        RECT 74.055 87.335 74.345 87.505 ;
        RECT 74.515 87.335 74.805 87.505 ;
        RECT 74.975 87.335 75.265 87.505 ;
        RECT 75.435 87.335 75.725 87.505 ;
        RECT 75.895 87.335 76.185 87.505 ;
        RECT 76.355 87.335 76.645 87.505 ;
        RECT 76.815 87.335 77.105 87.505 ;
        RECT 77.275 87.335 77.565 87.505 ;
        RECT 77.735 87.335 78.025 87.505 ;
        RECT 78.195 87.335 78.485 87.505 ;
        RECT 78.655 87.335 78.945 87.505 ;
        RECT 79.115 87.335 79.405 87.505 ;
        RECT 79.575 87.335 79.865 87.505 ;
        RECT 80.035 87.335 80.325 87.505 ;
        RECT 80.495 87.335 80.785 87.505 ;
        RECT 80.955 87.335 81.245 87.505 ;
        RECT 81.415 87.335 81.705 87.505 ;
        RECT 81.875 87.335 82.165 87.505 ;
        RECT 82.335 87.335 82.625 87.505 ;
        RECT 82.795 87.335 83.085 87.505 ;
        RECT 83.255 87.335 83.545 87.505 ;
        RECT 83.715 87.335 84.005 87.505 ;
        RECT 84.175 87.335 84.465 87.505 ;
        RECT 84.635 87.335 84.925 87.505 ;
        RECT 85.095 87.335 85.385 87.505 ;
        RECT 85.555 87.335 85.845 87.505 ;
        RECT 86.015 87.335 86.305 87.505 ;
        RECT 86.475 87.335 86.765 87.505 ;
        RECT 86.935 87.335 87.225 87.505 ;
        RECT 87.395 87.335 87.685 87.505 ;
        RECT 87.855 87.335 88.145 87.505 ;
        RECT 88.315 87.335 88.605 87.505 ;
        RECT 88.775 87.335 89.065 87.505 ;
        RECT 89.235 87.335 89.525 87.505 ;
        RECT 89.695 87.335 89.985 87.505 ;
        RECT 90.155 87.335 90.445 87.505 ;
        RECT 90.615 87.335 90.905 87.505 ;
        RECT 91.075 87.335 91.365 87.505 ;
        RECT 91.535 87.335 91.825 87.505 ;
        RECT 91.995 87.335 92.285 87.505 ;
        RECT 92.455 87.335 92.745 87.505 ;
        RECT 92.915 87.335 93.205 87.505 ;
        RECT 93.375 87.335 93.665 87.505 ;
        RECT 93.835 87.335 94.125 87.505 ;
        RECT 94.295 87.335 94.585 87.505 ;
        RECT 94.755 87.335 95.045 87.505 ;
        RECT 95.215 87.335 95.505 87.505 ;
        RECT 95.675 87.335 95.965 87.505 ;
        RECT 96.135 87.335 96.425 87.505 ;
        RECT 96.595 87.335 96.885 87.505 ;
        RECT 97.055 87.335 97.345 87.505 ;
        RECT 97.515 87.335 97.805 87.505 ;
        RECT 97.975 87.335 98.265 87.505 ;
        RECT 98.435 87.335 98.725 87.505 ;
        RECT 98.895 87.335 99.185 87.505 ;
        RECT 99.355 87.335 99.645 87.505 ;
        RECT 99.815 87.335 99.960 87.505 ;
        RECT 16.785 86.245 17.995 87.335 ;
        RECT 18.165 86.245 23.510 87.335 ;
        RECT 23.685 86.245 29.030 87.335 ;
        RECT 29.205 86.245 34.550 87.335 ;
        RECT 34.725 86.245 40.070 87.335 ;
        RECT 40.245 86.245 43.755 87.335 ;
        RECT 16.785 85.535 17.305 86.075 ;
        RECT 17.475 85.705 17.995 86.245 ;
        RECT 18.165 85.555 20.745 86.075 ;
        RECT 20.915 85.725 23.510 86.245 ;
        RECT 23.685 85.555 26.265 86.075 ;
        RECT 26.435 85.725 29.030 86.245 ;
        RECT 29.205 85.555 31.785 86.075 ;
        RECT 31.955 85.725 34.550 86.245 ;
        RECT 34.725 85.555 37.305 86.075 ;
        RECT 37.475 85.725 40.070 86.245 ;
        RECT 40.245 85.555 41.895 86.075 ;
        RECT 42.065 85.725 43.755 86.245 ;
        RECT 44.845 86.170 45.135 87.335 ;
        RECT 45.305 86.245 50.650 87.335 ;
        RECT 50.825 86.245 56.170 87.335 ;
        RECT 56.345 86.245 61.690 87.335 ;
        RECT 61.865 86.245 67.210 87.335 ;
        RECT 67.385 86.245 72.730 87.335 ;
        RECT 45.305 85.555 47.885 86.075 ;
        RECT 48.055 85.725 50.650 86.245 ;
        RECT 50.825 85.555 53.405 86.075 ;
        RECT 53.575 85.725 56.170 86.245 ;
        RECT 56.345 85.555 58.925 86.075 ;
        RECT 59.095 85.725 61.690 86.245 ;
        RECT 61.865 85.555 64.445 86.075 ;
        RECT 64.615 85.725 67.210 86.245 ;
        RECT 67.385 85.555 69.965 86.075 ;
        RECT 70.135 85.725 72.730 86.245 ;
        RECT 72.905 86.170 73.195 87.335 ;
        RECT 73.365 86.245 78.710 87.335 ;
        RECT 78.885 86.245 84.230 87.335 ;
        RECT 84.405 86.245 89.750 87.335 ;
        RECT 89.925 86.245 95.270 87.335 ;
        RECT 95.445 86.245 98.035 87.335 ;
        RECT 73.365 85.555 75.945 86.075 ;
        RECT 76.115 85.725 78.710 86.245 ;
        RECT 78.885 85.555 81.465 86.075 ;
        RECT 81.635 85.725 84.230 86.245 ;
        RECT 84.405 85.555 86.985 86.075 ;
        RECT 87.155 85.725 89.750 86.245 ;
        RECT 89.925 85.555 92.505 86.075 ;
        RECT 92.675 85.725 95.270 86.245 ;
        RECT 95.445 85.555 96.655 86.075 ;
        RECT 96.825 85.725 98.035 86.245 ;
        RECT 98.665 86.245 99.875 87.335 ;
        RECT 98.665 85.705 99.185 86.245 ;
        RECT 16.785 84.785 17.995 85.535 ;
        RECT 18.165 84.785 23.510 85.555 ;
        RECT 23.685 84.785 29.030 85.555 ;
        RECT 29.205 84.785 34.550 85.555 ;
        RECT 34.725 84.785 40.070 85.555 ;
        RECT 40.245 84.785 43.755 85.555 ;
        RECT 44.845 84.785 45.135 85.510 ;
        RECT 45.305 84.785 50.650 85.555 ;
        RECT 50.825 84.785 56.170 85.555 ;
        RECT 56.345 84.785 61.690 85.555 ;
        RECT 61.865 84.785 67.210 85.555 ;
        RECT 67.385 84.785 72.730 85.555 ;
        RECT 72.905 84.785 73.195 85.510 ;
        RECT 73.365 84.785 78.710 85.555 ;
        RECT 78.885 84.785 84.230 85.555 ;
        RECT 84.405 84.785 89.750 85.555 ;
        RECT 89.925 84.785 95.270 85.555 ;
        RECT 95.445 84.785 98.035 85.555 ;
        RECT 99.355 85.535 99.875 86.075 ;
        RECT 98.665 84.785 99.875 85.535 ;
        RECT 16.700 84.615 16.845 84.785 ;
        RECT 17.015 84.615 17.305 84.785 ;
        RECT 17.475 84.615 17.765 84.785 ;
        RECT 17.935 84.615 18.225 84.785 ;
        RECT 18.395 84.615 18.685 84.785 ;
        RECT 18.855 84.615 19.145 84.785 ;
        RECT 19.315 84.615 19.605 84.785 ;
        RECT 19.775 84.615 20.065 84.785 ;
        RECT 20.235 84.615 20.525 84.785 ;
        RECT 20.695 84.615 20.985 84.785 ;
        RECT 21.155 84.615 21.445 84.785 ;
        RECT 21.615 84.615 21.905 84.785 ;
        RECT 22.075 84.615 22.365 84.785 ;
        RECT 22.535 84.615 22.825 84.785 ;
        RECT 22.995 84.615 23.285 84.785 ;
        RECT 23.455 84.615 23.745 84.785 ;
        RECT 23.915 84.615 24.205 84.785 ;
        RECT 24.375 84.615 24.665 84.785 ;
        RECT 24.835 84.615 25.125 84.785 ;
        RECT 25.295 84.615 25.585 84.785 ;
        RECT 25.755 84.615 26.045 84.785 ;
        RECT 26.215 84.615 26.505 84.785 ;
        RECT 26.675 84.615 26.965 84.785 ;
        RECT 27.135 84.615 27.425 84.785 ;
        RECT 27.595 84.615 27.885 84.785 ;
        RECT 28.055 84.615 28.345 84.785 ;
        RECT 28.515 84.615 28.805 84.785 ;
        RECT 28.975 84.615 29.265 84.785 ;
        RECT 29.435 84.615 29.725 84.785 ;
        RECT 29.895 84.615 30.185 84.785 ;
        RECT 30.355 84.615 30.645 84.785 ;
        RECT 30.815 84.615 31.105 84.785 ;
        RECT 31.275 84.615 31.565 84.785 ;
        RECT 31.735 84.615 32.025 84.785 ;
        RECT 32.195 84.615 32.485 84.785 ;
        RECT 32.655 84.615 32.945 84.785 ;
        RECT 33.115 84.615 33.405 84.785 ;
        RECT 33.575 84.615 33.865 84.785 ;
        RECT 34.035 84.615 34.325 84.785 ;
        RECT 34.495 84.615 34.785 84.785 ;
        RECT 34.955 84.615 35.245 84.785 ;
        RECT 35.415 84.615 35.705 84.785 ;
        RECT 35.875 84.615 36.165 84.785 ;
        RECT 36.335 84.615 36.625 84.785 ;
        RECT 36.795 84.615 37.085 84.785 ;
        RECT 37.255 84.615 37.545 84.785 ;
        RECT 37.715 84.615 38.005 84.785 ;
        RECT 38.175 84.615 38.465 84.785 ;
        RECT 38.635 84.615 38.925 84.785 ;
        RECT 39.095 84.615 39.385 84.785 ;
        RECT 39.555 84.615 39.845 84.785 ;
        RECT 40.015 84.615 40.305 84.785 ;
        RECT 40.475 84.615 40.765 84.785 ;
        RECT 40.935 84.615 41.225 84.785 ;
        RECT 41.395 84.615 41.685 84.785 ;
        RECT 41.855 84.615 42.145 84.785 ;
        RECT 42.315 84.615 42.605 84.785 ;
        RECT 42.775 84.615 43.065 84.785 ;
        RECT 43.235 84.615 43.525 84.785 ;
        RECT 43.695 84.615 43.985 84.785 ;
        RECT 44.155 84.615 44.445 84.785 ;
        RECT 44.615 84.615 44.905 84.785 ;
        RECT 45.075 84.615 45.365 84.785 ;
        RECT 45.535 84.615 45.825 84.785 ;
        RECT 45.995 84.615 46.285 84.785 ;
        RECT 46.455 84.615 46.745 84.785 ;
        RECT 46.915 84.615 47.205 84.785 ;
        RECT 47.375 84.615 47.665 84.785 ;
        RECT 47.835 84.615 48.125 84.785 ;
        RECT 48.295 84.615 48.585 84.785 ;
        RECT 48.755 84.615 49.045 84.785 ;
        RECT 49.215 84.615 49.505 84.785 ;
        RECT 49.675 84.615 49.965 84.785 ;
        RECT 50.135 84.615 50.425 84.785 ;
        RECT 50.595 84.615 50.885 84.785 ;
        RECT 51.055 84.615 51.345 84.785 ;
        RECT 51.515 84.615 51.805 84.785 ;
        RECT 51.975 84.615 52.265 84.785 ;
        RECT 52.435 84.615 52.725 84.785 ;
        RECT 52.895 84.615 53.185 84.785 ;
        RECT 53.355 84.615 53.645 84.785 ;
        RECT 53.815 84.615 54.105 84.785 ;
        RECT 54.275 84.615 54.565 84.785 ;
        RECT 54.735 84.615 55.025 84.785 ;
        RECT 55.195 84.615 55.485 84.785 ;
        RECT 55.655 84.615 55.945 84.785 ;
        RECT 56.115 84.615 56.405 84.785 ;
        RECT 56.575 84.615 56.865 84.785 ;
        RECT 57.035 84.615 57.325 84.785 ;
        RECT 57.495 84.615 57.785 84.785 ;
        RECT 57.955 84.615 58.245 84.785 ;
        RECT 58.415 84.615 58.705 84.785 ;
        RECT 58.875 84.615 59.165 84.785 ;
        RECT 59.335 84.615 59.625 84.785 ;
        RECT 59.795 84.615 60.085 84.785 ;
        RECT 60.255 84.615 60.545 84.785 ;
        RECT 60.715 84.615 61.005 84.785 ;
        RECT 61.175 84.615 61.465 84.785 ;
        RECT 61.635 84.615 61.925 84.785 ;
        RECT 62.095 84.615 62.385 84.785 ;
        RECT 62.555 84.615 62.845 84.785 ;
        RECT 63.015 84.615 63.305 84.785 ;
        RECT 63.475 84.615 63.765 84.785 ;
        RECT 63.935 84.615 64.225 84.785 ;
        RECT 64.395 84.615 64.685 84.785 ;
        RECT 64.855 84.615 65.145 84.785 ;
        RECT 65.315 84.615 65.605 84.785 ;
        RECT 65.775 84.615 66.065 84.785 ;
        RECT 66.235 84.615 66.525 84.785 ;
        RECT 66.695 84.615 66.985 84.785 ;
        RECT 67.155 84.615 67.445 84.785 ;
        RECT 67.615 84.615 67.905 84.785 ;
        RECT 68.075 84.615 68.365 84.785 ;
        RECT 68.535 84.615 68.825 84.785 ;
        RECT 68.995 84.615 69.285 84.785 ;
        RECT 69.455 84.615 69.745 84.785 ;
        RECT 69.915 84.615 70.205 84.785 ;
        RECT 70.375 84.615 70.665 84.785 ;
        RECT 70.835 84.615 71.125 84.785 ;
        RECT 71.295 84.615 71.585 84.785 ;
        RECT 71.755 84.615 72.045 84.785 ;
        RECT 72.215 84.615 72.505 84.785 ;
        RECT 72.675 84.615 72.965 84.785 ;
        RECT 73.135 84.615 73.425 84.785 ;
        RECT 73.595 84.615 73.885 84.785 ;
        RECT 74.055 84.615 74.345 84.785 ;
        RECT 74.515 84.615 74.805 84.785 ;
        RECT 74.975 84.615 75.265 84.785 ;
        RECT 75.435 84.615 75.725 84.785 ;
        RECT 75.895 84.615 76.185 84.785 ;
        RECT 76.355 84.615 76.645 84.785 ;
        RECT 76.815 84.615 77.105 84.785 ;
        RECT 77.275 84.615 77.565 84.785 ;
        RECT 77.735 84.615 78.025 84.785 ;
        RECT 78.195 84.615 78.485 84.785 ;
        RECT 78.655 84.615 78.945 84.785 ;
        RECT 79.115 84.615 79.405 84.785 ;
        RECT 79.575 84.615 79.865 84.785 ;
        RECT 80.035 84.615 80.325 84.785 ;
        RECT 80.495 84.615 80.785 84.785 ;
        RECT 80.955 84.615 81.245 84.785 ;
        RECT 81.415 84.615 81.705 84.785 ;
        RECT 81.875 84.615 82.165 84.785 ;
        RECT 82.335 84.615 82.625 84.785 ;
        RECT 82.795 84.615 83.085 84.785 ;
        RECT 83.255 84.615 83.545 84.785 ;
        RECT 83.715 84.615 84.005 84.785 ;
        RECT 84.175 84.615 84.465 84.785 ;
        RECT 84.635 84.615 84.925 84.785 ;
        RECT 85.095 84.615 85.385 84.785 ;
        RECT 85.555 84.615 85.845 84.785 ;
        RECT 86.015 84.615 86.305 84.785 ;
        RECT 86.475 84.615 86.765 84.785 ;
        RECT 86.935 84.615 87.225 84.785 ;
        RECT 87.395 84.615 87.685 84.785 ;
        RECT 87.855 84.615 88.145 84.785 ;
        RECT 88.315 84.615 88.605 84.785 ;
        RECT 88.775 84.615 89.065 84.785 ;
        RECT 89.235 84.615 89.525 84.785 ;
        RECT 89.695 84.615 89.985 84.785 ;
        RECT 90.155 84.615 90.445 84.785 ;
        RECT 90.615 84.615 90.905 84.785 ;
        RECT 91.075 84.615 91.365 84.785 ;
        RECT 91.535 84.615 91.825 84.785 ;
        RECT 91.995 84.615 92.285 84.785 ;
        RECT 92.455 84.615 92.745 84.785 ;
        RECT 92.915 84.615 93.205 84.785 ;
        RECT 93.375 84.615 93.665 84.785 ;
        RECT 93.835 84.615 94.125 84.785 ;
        RECT 94.295 84.615 94.585 84.785 ;
        RECT 94.755 84.615 95.045 84.785 ;
        RECT 95.215 84.615 95.505 84.785 ;
        RECT 95.675 84.615 95.965 84.785 ;
        RECT 96.135 84.615 96.425 84.785 ;
        RECT 96.595 84.615 96.885 84.785 ;
        RECT 97.055 84.615 97.345 84.785 ;
        RECT 97.515 84.615 97.805 84.785 ;
        RECT 97.975 84.615 98.265 84.785 ;
        RECT 98.435 84.615 98.725 84.785 ;
        RECT 98.895 84.615 99.185 84.785 ;
        RECT 99.355 84.615 99.645 84.785 ;
        RECT 99.815 84.615 99.960 84.785 ;
        RECT 16.785 83.865 17.995 84.615 ;
        RECT 16.785 83.325 17.305 83.865 ;
        RECT 18.165 83.845 23.510 84.615 ;
        RECT 23.685 83.845 29.030 84.615 ;
        RECT 29.205 83.845 30.875 84.615 ;
        RECT 31.045 83.890 31.335 84.615 ;
        RECT 31.505 83.845 35.015 84.615 ;
        RECT 17.475 83.155 17.995 83.695 ;
        RECT 18.165 83.325 20.745 83.845 ;
        RECT 20.915 83.155 23.510 83.675 ;
        RECT 23.685 83.325 26.265 83.845 ;
        RECT 26.435 83.155 29.030 83.675 ;
        RECT 29.205 83.325 29.955 83.845 ;
        RECT 30.125 83.155 30.875 83.675 ;
        RECT 31.505 83.325 33.155 83.845 ;
        RECT 35.225 83.795 35.455 84.615 ;
      LAYER li1 ;
        RECT 35.625 83.815 35.955 84.445 ;
      LAYER li1 ;
        RECT 16.785 82.065 17.995 83.155 ;
        RECT 18.165 82.065 23.510 83.155 ;
        RECT 23.685 82.065 29.030 83.155 ;
        RECT 29.205 82.065 30.875 83.155 ;
        RECT 31.045 82.065 31.335 83.230 ;
        RECT 33.325 83.155 35.015 83.675 ;
      LAYER li1 ;
        RECT 35.705 83.215 35.955 83.815 ;
      LAYER li1 ;
        RECT 36.125 83.795 36.335 84.615 ;
        RECT 36.565 83.845 41.910 84.615 ;
        RECT 42.085 83.845 47.430 84.615 ;
        RECT 47.605 83.845 52.950 84.615 ;
        RECT 53.125 83.845 58.470 84.615 ;
        RECT 59.105 83.890 59.395 84.615 ;
        RECT 59.565 83.845 64.910 84.615 ;
        RECT 65.085 83.845 70.430 84.615 ;
        RECT 70.605 83.845 75.950 84.615 ;
        RECT 76.125 83.845 81.470 84.615 ;
        RECT 81.645 83.845 86.990 84.615 ;
        RECT 87.165 83.890 87.455 84.615 ;
        RECT 87.625 83.845 92.970 84.615 ;
        RECT 93.145 83.845 98.490 84.615 ;
        RECT 98.665 83.865 99.875 84.615 ;
        RECT 36.565 83.325 39.145 83.845 ;
        RECT 31.505 82.065 35.015 83.155 ;
        RECT 35.225 82.065 35.455 83.205 ;
      LAYER li1 ;
        RECT 35.625 82.235 35.955 83.215 ;
      LAYER li1 ;
        RECT 36.125 82.065 36.335 83.205 ;
        RECT 39.315 83.155 41.910 83.675 ;
        RECT 42.085 83.325 44.665 83.845 ;
        RECT 44.835 83.155 47.430 83.675 ;
        RECT 47.605 83.325 50.185 83.845 ;
        RECT 50.355 83.155 52.950 83.675 ;
        RECT 53.125 83.325 55.705 83.845 ;
        RECT 55.875 83.155 58.470 83.675 ;
        RECT 59.565 83.325 62.145 83.845 ;
        RECT 36.565 82.065 41.910 83.155 ;
        RECT 42.085 82.065 47.430 83.155 ;
        RECT 47.605 82.065 52.950 83.155 ;
        RECT 53.125 82.065 58.470 83.155 ;
        RECT 59.105 82.065 59.395 83.230 ;
        RECT 62.315 83.155 64.910 83.675 ;
        RECT 65.085 83.325 67.665 83.845 ;
        RECT 67.835 83.155 70.430 83.675 ;
        RECT 70.605 83.325 73.185 83.845 ;
        RECT 73.355 83.155 75.950 83.675 ;
        RECT 76.125 83.325 78.705 83.845 ;
        RECT 78.875 83.155 81.470 83.675 ;
        RECT 81.645 83.325 84.225 83.845 ;
        RECT 84.395 83.155 86.990 83.675 ;
        RECT 87.625 83.325 90.205 83.845 ;
        RECT 59.565 82.065 64.910 83.155 ;
        RECT 65.085 82.065 70.430 83.155 ;
        RECT 70.605 82.065 75.950 83.155 ;
        RECT 76.125 82.065 81.470 83.155 ;
        RECT 81.645 82.065 86.990 83.155 ;
        RECT 87.165 82.065 87.455 83.230 ;
        RECT 90.375 83.155 92.970 83.675 ;
        RECT 93.145 83.325 95.725 83.845 ;
        RECT 95.895 83.155 98.490 83.675 ;
        RECT 87.625 82.065 92.970 83.155 ;
        RECT 93.145 82.065 98.490 83.155 ;
        RECT 98.665 83.155 99.185 83.695 ;
        RECT 99.355 83.325 99.875 83.865 ;
        RECT 98.665 82.065 99.875 83.155 ;
        RECT 16.700 81.895 16.845 82.065 ;
        RECT 17.015 81.895 17.305 82.065 ;
        RECT 17.475 81.895 17.765 82.065 ;
        RECT 17.935 81.895 18.225 82.065 ;
        RECT 18.395 81.895 18.685 82.065 ;
        RECT 18.855 81.895 19.145 82.065 ;
        RECT 19.315 81.895 19.605 82.065 ;
        RECT 19.775 81.895 20.065 82.065 ;
        RECT 20.235 81.895 20.525 82.065 ;
        RECT 20.695 81.895 20.985 82.065 ;
        RECT 21.155 81.895 21.445 82.065 ;
        RECT 21.615 81.895 21.905 82.065 ;
        RECT 22.075 81.895 22.365 82.065 ;
        RECT 22.535 81.895 22.825 82.065 ;
        RECT 22.995 81.895 23.285 82.065 ;
        RECT 23.455 81.895 23.745 82.065 ;
        RECT 23.915 81.895 24.205 82.065 ;
        RECT 24.375 81.895 24.665 82.065 ;
        RECT 24.835 81.895 25.125 82.065 ;
        RECT 25.295 81.895 25.585 82.065 ;
        RECT 25.755 81.895 26.045 82.065 ;
        RECT 26.215 81.895 26.505 82.065 ;
        RECT 26.675 81.895 26.965 82.065 ;
        RECT 27.135 81.895 27.425 82.065 ;
        RECT 27.595 81.895 27.885 82.065 ;
        RECT 28.055 81.895 28.345 82.065 ;
        RECT 28.515 81.895 28.805 82.065 ;
        RECT 28.975 81.895 29.265 82.065 ;
        RECT 29.435 81.895 29.725 82.065 ;
        RECT 29.895 81.895 30.185 82.065 ;
        RECT 30.355 81.895 30.645 82.065 ;
        RECT 30.815 81.895 31.105 82.065 ;
        RECT 31.275 81.895 31.565 82.065 ;
        RECT 31.735 81.895 32.025 82.065 ;
        RECT 32.195 81.895 32.485 82.065 ;
        RECT 32.655 81.895 32.945 82.065 ;
        RECT 33.115 81.895 33.405 82.065 ;
        RECT 33.575 81.895 33.865 82.065 ;
        RECT 34.035 81.895 34.325 82.065 ;
        RECT 34.495 81.895 34.785 82.065 ;
        RECT 34.955 81.895 35.245 82.065 ;
        RECT 35.415 81.895 35.705 82.065 ;
        RECT 35.875 81.895 36.165 82.065 ;
        RECT 36.335 81.895 36.625 82.065 ;
        RECT 36.795 81.895 37.085 82.065 ;
        RECT 37.255 81.895 37.545 82.065 ;
        RECT 37.715 81.895 38.005 82.065 ;
        RECT 38.175 81.895 38.465 82.065 ;
        RECT 38.635 81.895 38.925 82.065 ;
        RECT 39.095 81.895 39.385 82.065 ;
        RECT 39.555 81.895 39.845 82.065 ;
        RECT 40.015 81.895 40.305 82.065 ;
        RECT 40.475 81.895 40.765 82.065 ;
        RECT 40.935 81.895 41.225 82.065 ;
        RECT 41.395 81.895 41.685 82.065 ;
        RECT 41.855 81.895 42.145 82.065 ;
        RECT 42.315 81.895 42.605 82.065 ;
        RECT 42.775 81.895 43.065 82.065 ;
        RECT 43.235 81.895 43.525 82.065 ;
        RECT 43.695 81.895 43.985 82.065 ;
        RECT 44.155 81.895 44.445 82.065 ;
        RECT 44.615 81.895 44.905 82.065 ;
        RECT 45.075 81.895 45.365 82.065 ;
        RECT 45.535 81.895 45.825 82.065 ;
        RECT 45.995 81.895 46.285 82.065 ;
        RECT 46.455 81.895 46.745 82.065 ;
        RECT 46.915 81.895 47.205 82.065 ;
        RECT 47.375 81.895 47.665 82.065 ;
        RECT 47.835 81.895 48.125 82.065 ;
        RECT 48.295 81.895 48.585 82.065 ;
        RECT 48.755 81.895 49.045 82.065 ;
        RECT 49.215 81.895 49.505 82.065 ;
        RECT 49.675 81.895 49.965 82.065 ;
        RECT 50.135 81.895 50.425 82.065 ;
        RECT 50.595 81.895 50.885 82.065 ;
        RECT 51.055 81.895 51.345 82.065 ;
        RECT 51.515 81.895 51.805 82.065 ;
        RECT 51.975 81.895 52.265 82.065 ;
        RECT 52.435 81.895 52.725 82.065 ;
        RECT 52.895 81.895 53.185 82.065 ;
        RECT 53.355 81.895 53.645 82.065 ;
        RECT 53.815 81.895 54.105 82.065 ;
        RECT 54.275 81.895 54.565 82.065 ;
        RECT 54.735 81.895 55.025 82.065 ;
        RECT 55.195 81.895 55.485 82.065 ;
        RECT 55.655 81.895 55.945 82.065 ;
        RECT 56.115 81.895 56.405 82.065 ;
        RECT 56.575 81.895 56.865 82.065 ;
        RECT 57.035 81.895 57.325 82.065 ;
        RECT 57.495 81.895 57.785 82.065 ;
        RECT 57.955 81.895 58.245 82.065 ;
        RECT 58.415 81.895 58.705 82.065 ;
        RECT 58.875 81.895 59.165 82.065 ;
        RECT 59.335 81.895 59.625 82.065 ;
        RECT 59.795 81.895 60.085 82.065 ;
        RECT 60.255 81.895 60.545 82.065 ;
        RECT 60.715 81.895 61.005 82.065 ;
        RECT 61.175 81.895 61.465 82.065 ;
        RECT 61.635 81.895 61.925 82.065 ;
        RECT 62.095 81.895 62.385 82.065 ;
        RECT 62.555 81.895 62.845 82.065 ;
        RECT 63.015 81.895 63.305 82.065 ;
        RECT 63.475 81.895 63.765 82.065 ;
        RECT 63.935 81.895 64.225 82.065 ;
        RECT 64.395 81.895 64.685 82.065 ;
        RECT 64.855 81.895 65.145 82.065 ;
        RECT 65.315 81.895 65.605 82.065 ;
        RECT 65.775 81.895 66.065 82.065 ;
        RECT 66.235 81.895 66.525 82.065 ;
        RECT 66.695 81.895 66.985 82.065 ;
        RECT 67.155 81.895 67.445 82.065 ;
        RECT 67.615 81.895 67.905 82.065 ;
        RECT 68.075 81.895 68.365 82.065 ;
        RECT 68.535 81.895 68.825 82.065 ;
        RECT 68.995 81.895 69.285 82.065 ;
        RECT 69.455 81.895 69.745 82.065 ;
        RECT 69.915 81.895 70.205 82.065 ;
        RECT 70.375 81.895 70.665 82.065 ;
        RECT 70.835 81.895 71.125 82.065 ;
        RECT 71.295 81.895 71.585 82.065 ;
        RECT 71.755 81.895 72.045 82.065 ;
        RECT 72.215 81.895 72.505 82.065 ;
        RECT 72.675 81.895 72.965 82.065 ;
        RECT 73.135 81.895 73.425 82.065 ;
        RECT 73.595 81.895 73.885 82.065 ;
        RECT 74.055 81.895 74.345 82.065 ;
        RECT 74.515 81.895 74.805 82.065 ;
        RECT 74.975 81.895 75.265 82.065 ;
        RECT 75.435 81.895 75.725 82.065 ;
        RECT 75.895 81.895 76.185 82.065 ;
        RECT 76.355 81.895 76.645 82.065 ;
        RECT 76.815 81.895 77.105 82.065 ;
        RECT 77.275 81.895 77.565 82.065 ;
        RECT 77.735 81.895 78.025 82.065 ;
        RECT 78.195 81.895 78.485 82.065 ;
        RECT 78.655 81.895 78.945 82.065 ;
        RECT 79.115 81.895 79.405 82.065 ;
        RECT 79.575 81.895 79.865 82.065 ;
        RECT 80.035 81.895 80.325 82.065 ;
        RECT 80.495 81.895 80.785 82.065 ;
        RECT 80.955 81.895 81.245 82.065 ;
        RECT 81.415 81.895 81.705 82.065 ;
        RECT 81.875 81.895 82.165 82.065 ;
        RECT 82.335 81.895 82.625 82.065 ;
        RECT 82.795 81.895 83.085 82.065 ;
        RECT 83.255 81.895 83.545 82.065 ;
        RECT 83.715 81.895 84.005 82.065 ;
        RECT 84.175 81.895 84.465 82.065 ;
        RECT 84.635 81.895 84.925 82.065 ;
        RECT 85.095 81.895 85.385 82.065 ;
        RECT 85.555 81.895 85.845 82.065 ;
        RECT 86.015 81.895 86.305 82.065 ;
        RECT 86.475 81.895 86.765 82.065 ;
        RECT 86.935 81.895 87.225 82.065 ;
        RECT 87.395 81.895 87.685 82.065 ;
        RECT 87.855 81.895 88.145 82.065 ;
        RECT 88.315 81.895 88.605 82.065 ;
        RECT 88.775 81.895 89.065 82.065 ;
        RECT 89.235 81.895 89.525 82.065 ;
        RECT 89.695 81.895 89.985 82.065 ;
        RECT 90.155 81.895 90.445 82.065 ;
        RECT 90.615 81.895 90.905 82.065 ;
        RECT 91.075 81.895 91.365 82.065 ;
        RECT 91.535 81.895 91.825 82.065 ;
        RECT 91.995 81.895 92.285 82.065 ;
        RECT 92.455 81.895 92.745 82.065 ;
        RECT 92.915 81.895 93.205 82.065 ;
        RECT 93.375 81.895 93.665 82.065 ;
        RECT 93.835 81.895 94.125 82.065 ;
        RECT 94.295 81.895 94.585 82.065 ;
        RECT 94.755 81.895 95.045 82.065 ;
        RECT 95.215 81.895 95.505 82.065 ;
        RECT 95.675 81.895 95.965 82.065 ;
        RECT 96.135 81.895 96.425 82.065 ;
        RECT 96.595 81.895 96.885 82.065 ;
        RECT 97.055 81.895 97.345 82.065 ;
        RECT 97.515 81.895 97.805 82.065 ;
        RECT 97.975 81.895 98.265 82.065 ;
        RECT 98.435 81.895 98.725 82.065 ;
        RECT 98.895 81.895 99.185 82.065 ;
        RECT 99.355 81.895 99.645 82.065 ;
        RECT 99.815 81.895 99.960 82.065 ;
        RECT 16.785 80.805 17.995 81.895 ;
        RECT 18.165 80.805 23.510 81.895 ;
        RECT 23.685 80.805 29.030 81.895 ;
        RECT 29.205 80.805 34.550 81.895 ;
        RECT 34.725 80.805 37.315 81.895 ;
        RECT 37.955 81.140 38.285 81.895 ;
        RECT 38.465 81.010 38.645 81.725 ;
        RECT 38.850 81.195 39.180 81.895 ;
      LAYER li1 ;
        RECT 39.390 81.020 39.580 81.725 ;
      LAYER li1 ;
        RECT 39.750 81.195 40.080 81.895 ;
      LAYER li1 ;
        RECT 40.250 81.025 40.440 81.725 ;
      LAYER li1 ;
        RECT 40.610 81.195 40.940 81.895 ;
      LAYER li1 ;
        RECT 40.250 81.020 40.995 81.025 ;
      LAYER li1 ;
        RECT 16.785 80.095 17.305 80.635 ;
        RECT 17.475 80.265 17.995 80.805 ;
        RECT 18.165 80.115 20.745 80.635 ;
        RECT 20.915 80.285 23.510 80.805 ;
        RECT 23.685 80.115 26.265 80.635 ;
        RECT 26.435 80.285 29.030 80.805 ;
        RECT 29.205 80.115 31.785 80.635 ;
        RECT 31.955 80.285 34.550 80.805 ;
        RECT 34.725 80.115 35.935 80.635 ;
        RECT 36.105 80.285 37.315 80.805 ;
      LAYER li1 ;
        RECT 37.985 80.255 38.295 80.875 ;
      LAYER li1 ;
        RECT 38.465 80.840 39.220 81.010 ;
        RECT 39.010 80.615 39.220 80.840 ;
      LAYER li1 ;
        RECT 39.390 80.795 40.995 81.020 ;
      LAYER li1 ;
        RECT 41.165 80.805 44.675 81.895 ;
        RECT 39.010 80.280 40.545 80.615 ;
        RECT 16.785 79.345 17.995 80.095 ;
        RECT 18.165 79.345 23.510 80.115 ;
        RECT 23.685 79.345 29.030 80.115 ;
        RECT 29.205 79.345 34.550 80.115 ;
        RECT 34.725 79.345 37.315 80.115 ;
        RECT 39.010 80.065 39.220 80.280 ;
      LAYER li1 ;
        RECT 40.715 80.105 40.995 80.795 ;
      LAYER li1 ;
        RECT 37.955 79.875 39.220 80.065 ;
      LAYER li1 ;
        RECT 39.390 79.875 40.995 80.105 ;
      LAYER li1 ;
        RECT 41.165 80.115 42.815 80.635 ;
        RECT 42.985 80.285 44.675 80.805 ;
        RECT 44.845 80.730 45.135 81.895 ;
        RECT 45.305 80.805 50.650 81.895 ;
        RECT 50.825 80.805 56.170 81.895 ;
        RECT 56.345 80.805 61.690 81.895 ;
        RECT 61.865 80.805 67.210 81.895 ;
        RECT 67.385 80.805 72.730 81.895 ;
        RECT 45.305 80.115 47.885 80.635 ;
        RECT 48.055 80.285 50.650 80.805 ;
        RECT 50.825 80.115 53.405 80.635 ;
        RECT 53.575 80.285 56.170 80.805 ;
        RECT 56.345 80.115 58.925 80.635 ;
        RECT 59.095 80.285 61.690 80.805 ;
        RECT 61.865 80.115 64.445 80.635 ;
        RECT 64.615 80.285 67.210 80.805 ;
        RECT 67.385 80.115 69.965 80.635 ;
        RECT 70.135 80.285 72.730 80.805 ;
        RECT 72.905 80.730 73.195 81.895 ;
        RECT 73.365 80.805 78.710 81.895 ;
        RECT 78.885 80.805 84.230 81.895 ;
        RECT 84.405 80.805 89.750 81.895 ;
        RECT 89.925 80.805 95.270 81.895 ;
        RECT 95.445 80.805 98.035 81.895 ;
        RECT 73.365 80.115 75.945 80.635 ;
        RECT 76.115 80.285 78.710 80.805 ;
        RECT 78.885 80.115 81.465 80.635 ;
        RECT 81.635 80.285 84.230 80.805 ;
        RECT 84.405 80.115 86.985 80.635 ;
        RECT 87.155 80.285 89.750 80.805 ;
        RECT 89.925 80.115 92.505 80.635 ;
        RECT 92.675 80.285 95.270 80.805 ;
        RECT 95.445 80.115 96.655 80.635 ;
        RECT 96.825 80.285 98.035 80.805 ;
        RECT 98.665 80.805 99.875 81.895 ;
        RECT 98.665 80.265 99.185 80.805 ;
        RECT 37.955 79.515 38.285 79.875 ;
      LAYER li1 ;
        RECT 39.390 79.775 39.580 79.875 ;
      LAYER li1 ;
        RECT 38.815 79.345 39.145 79.705 ;
        RECT 39.750 79.345 40.080 79.705 ;
      LAYER li1 ;
        RECT 40.250 79.515 40.440 79.875 ;
      LAYER li1 ;
        RECT 40.610 79.345 40.940 79.705 ;
        RECT 41.165 79.345 44.675 80.115 ;
        RECT 44.845 79.345 45.135 80.070 ;
        RECT 45.305 79.345 50.650 80.115 ;
        RECT 50.825 79.345 56.170 80.115 ;
        RECT 56.345 79.345 61.690 80.115 ;
        RECT 61.865 79.345 67.210 80.115 ;
        RECT 67.385 79.345 72.730 80.115 ;
        RECT 72.905 79.345 73.195 80.070 ;
        RECT 73.365 79.345 78.710 80.115 ;
        RECT 78.885 79.345 84.230 80.115 ;
        RECT 84.405 79.345 89.750 80.115 ;
        RECT 89.925 79.345 95.270 80.115 ;
        RECT 95.445 79.345 98.035 80.115 ;
        RECT 99.355 80.095 99.875 80.635 ;
        RECT 98.665 79.345 99.875 80.095 ;
        RECT 16.700 79.175 16.845 79.345 ;
        RECT 17.015 79.175 17.305 79.345 ;
        RECT 17.475 79.175 17.765 79.345 ;
        RECT 17.935 79.175 18.225 79.345 ;
        RECT 18.395 79.175 18.685 79.345 ;
        RECT 18.855 79.175 19.145 79.345 ;
        RECT 19.315 79.175 19.605 79.345 ;
        RECT 19.775 79.175 20.065 79.345 ;
        RECT 20.235 79.175 20.525 79.345 ;
        RECT 20.695 79.175 20.985 79.345 ;
        RECT 21.155 79.175 21.445 79.345 ;
        RECT 21.615 79.175 21.905 79.345 ;
        RECT 22.075 79.175 22.365 79.345 ;
        RECT 22.535 79.175 22.825 79.345 ;
        RECT 22.995 79.175 23.285 79.345 ;
        RECT 23.455 79.175 23.745 79.345 ;
        RECT 23.915 79.175 24.205 79.345 ;
        RECT 24.375 79.175 24.665 79.345 ;
        RECT 24.835 79.175 25.125 79.345 ;
        RECT 25.295 79.175 25.585 79.345 ;
        RECT 25.755 79.175 26.045 79.345 ;
        RECT 26.215 79.175 26.505 79.345 ;
        RECT 26.675 79.175 26.965 79.345 ;
        RECT 27.135 79.175 27.425 79.345 ;
        RECT 27.595 79.175 27.885 79.345 ;
        RECT 28.055 79.175 28.345 79.345 ;
        RECT 28.515 79.175 28.805 79.345 ;
        RECT 28.975 79.175 29.265 79.345 ;
        RECT 29.435 79.175 29.725 79.345 ;
        RECT 29.895 79.175 30.185 79.345 ;
        RECT 30.355 79.175 30.645 79.345 ;
        RECT 30.815 79.175 31.105 79.345 ;
        RECT 31.275 79.175 31.565 79.345 ;
        RECT 31.735 79.175 32.025 79.345 ;
        RECT 32.195 79.175 32.485 79.345 ;
        RECT 32.655 79.175 32.945 79.345 ;
        RECT 33.115 79.175 33.405 79.345 ;
        RECT 33.575 79.175 33.865 79.345 ;
        RECT 34.035 79.175 34.325 79.345 ;
        RECT 34.495 79.175 34.785 79.345 ;
        RECT 34.955 79.175 35.245 79.345 ;
        RECT 35.415 79.175 35.705 79.345 ;
        RECT 35.875 79.175 36.165 79.345 ;
        RECT 36.335 79.175 36.625 79.345 ;
        RECT 36.795 79.175 37.085 79.345 ;
        RECT 37.255 79.175 37.545 79.345 ;
        RECT 37.715 79.175 38.005 79.345 ;
        RECT 38.175 79.175 38.465 79.345 ;
        RECT 38.635 79.175 38.925 79.345 ;
        RECT 39.095 79.175 39.385 79.345 ;
        RECT 39.555 79.175 39.845 79.345 ;
        RECT 40.015 79.175 40.305 79.345 ;
        RECT 40.475 79.175 40.765 79.345 ;
        RECT 40.935 79.175 41.225 79.345 ;
        RECT 41.395 79.175 41.685 79.345 ;
        RECT 41.855 79.175 42.145 79.345 ;
        RECT 42.315 79.175 42.605 79.345 ;
        RECT 42.775 79.175 43.065 79.345 ;
        RECT 43.235 79.175 43.525 79.345 ;
        RECT 43.695 79.175 43.985 79.345 ;
        RECT 44.155 79.175 44.445 79.345 ;
        RECT 44.615 79.175 44.905 79.345 ;
        RECT 45.075 79.175 45.365 79.345 ;
        RECT 45.535 79.175 45.825 79.345 ;
        RECT 45.995 79.175 46.285 79.345 ;
        RECT 46.455 79.175 46.745 79.345 ;
        RECT 46.915 79.175 47.205 79.345 ;
        RECT 47.375 79.175 47.665 79.345 ;
        RECT 47.835 79.175 48.125 79.345 ;
        RECT 48.295 79.175 48.585 79.345 ;
        RECT 48.755 79.175 49.045 79.345 ;
        RECT 49.215 79.175 49.505 79.345 ;
        RECT 49.675 79.175 49.965 79.345 ;
        RECT 50.135 79.175 50.425 79.345 ;
        RECT 50.595 79.175 50.885 79.345 ;
        RECT 51.055 79.175 51.345 79.345 ;
        RECT 51.515 79.175 51.805 79.345 ;
        RECT 51.975 79.175 52.265 79.345 ;
        RECT 52.435 79.175 52.725 79.345 ;
        RECT 52.895 79.175 53.185 79.345 ;
        RECT 53.355 79.175 53.645 79.345 ;
        RECT 53.815 79.175 54.105 79.345 ;
        RECT 54.275 79.175 54.565 79.345 ;
        RECT 54.735 79.175 55.025 79.345 ;
        RECT 55.195 79.175 55.485 79.345 ;
        RECT 55.655 79.175 55.945 79.345 ;
        RECT 56.115 79.175 56.405 79.345 ;
        RECT 56.575 79.175 56.865 79.345 ;
        RECT 57.035 79.175 57.325 79.345 ;
        RECT 57.495 79.175 57.785 79.345 ;
        RECT 57.955 79.175 58.245 79.345 ;
        RECT 58.415 79.175 58.705 79.345 ;
        RECT 58.875 79.175 59.165 79.345 ;
        RECT 59.335 79.175 59.625 79.345 ;
        RECT 59.795 79.175 60.085 79.345 ;
        RECT 60.255 79.175 60.545 79.345 ;
        RECT 60.715 79.175 61.005 79.345 ;
        RECT 61.175 79.175 61.465 79.345 ;
        RECT 61.635 79.175 61.925 79.345 ;
        RECT 62.095 79.175 62.385 79.345 ;
        RECT 62.555 79.175 62.845 79.345 ;
        RECT 63.015 79.175 63.305 79.345 ;
        RECT 63.475 79.175 63.765 79.345 ;
        RECT 63.935 79.175 64.225 79.345 ;
        RECT 64.395 79.175 64.685 79.345 ;
        RECT 64.855 79.175 65.145 79.345 ;
        RECT 65.315 79.175 65.605 79.345 ;
        RECT 65.775 79.175 66.065 79.345 ;
        RECT 66.235 79.175 66.525 79.345 ;
        RECT 66.695 79.175 66.985 79.345 ;
        RECT 67.155 79.175 67.445 79.345 ;
        RECT 67.615 79.175 67.905 79.345 ;
        RECT 68.075 79.175 68.365 79.345 ;
        RECT 68.535 79.175 68.825 79.345 ;
        RECT 68.995 79.175 69.285 79.345 ;
        RECT 69.455 79.175 69.745 79.345 ;
        RECT 69.915 79.175 70.205 79.345 ;
        RECT 70.375 79.175 70.665 79.345 ;
        RECT 70.835 79.175 71.125 79.345 ;
        RECT 71.295 79.175 71.585 79.345 ;
        RECT 71.755 79.175 72.045 79.345 ;
        RECT 72.215 79.175 72.505 79.345 ;
        RECT 72.675 79.175 72.965 79.345 ;
        RECT 73.135 79.175 73.425 79.345 ;
        RECT 73.595 79.175 73.885 79.345 ;
        RECT 74.055 79.175 74.345 79.345 ;
        RECT 74.515 79.175 74.805 79.345 ;
        RECT 74.975 79.175 75.265 79.345 ;
        RECT 75.435 79.175 75.725 79.345 ;
        RECT 75.895 79.175 76.185 79.345 ;
        RECT 76.355 79.175 76.645 79.345 ;
        RECT 76.815 79.175 77.105 79.345 ;
        RECT 77.275 79.175 77.565 79.345 ;
        RECT 77.735 79.175 78.025 79.345 ;
        RECT 78.195 79.175 78.485 79.345 ;
        RECT 78.655 79.175 78.945 79.345 ;
        RECT 79.115 79.175 79.405 79.345 ;
        RECT 79.575 79.175 79.865 79.345 ;
        RECT 80.035 79.175 80.325 79.345 ;
        RECT 80.495 79.175 80.785 79.345 ;
        RECT 80.955 79.175 81.245 79.345 ;
        RECT 81.415 79.175 81.705 79.345 ;
        RECT 81.875 79.175 82.165 79.345 ;
        RECT 82.335 79.175 82.625 79.345 ;
        RECT 82.795 79.175 83.085 79.345 ;
        RECT 83.255 79.175 83.545 79.345 ;
        RECT 83.715 79.175 84.005 79.345 ;
        RECT 84.175 79.175 84.465 79.345 ;
        RECT 84.635 79.175 84.925 79.345 ;
        RECT 85.095 79.175 85.385 79.345 ;
        RECT 85.555 79.175 85.845 79.345 ;
        RECT 86.015 79.175 86.305 79.345 ;
        RECT 86.475 79.175 86.765 79.345 ;
        RECT 86.935 79.175 87.225 79.345 ;
        RECT 87.395 79.175 87.685 79.345 ;
        RECT 87.855 79.175 88.145 79.345 ;
        RECT 88.315 79.175 88.605 79.345 ;
        RECT 88.775 79.175 89.065 79.345 ;
        RECT 89.235 79.175 89.525 79.345 ;
        RECT 89.695 79.175 89.985 79.345 ;
        RECT 90.155 79.175 90.445 79.345 ;
        RECT 90.615 79.175 90.905 79.345 ;
        RECT 91.075 79.175 91.365 79.345 ;
        RECT 91.535 79.175 91.825 79.345 ;
        RECT 91.995 79.175 92.285 79.345 ;
        RECT 92.455 79.175 92.745 79.345 ;
        RECT 92.915 79.175 93.205 79.345 ;
        RECT 93.375 79.175 93.665 79.345 ;
        RECT 93.835 79.175 94.125 79.345 ;
        RECT 94.295 79.175 94.585 79.345 ;
        RECT 94.755 79.175 95.045 79.345 ;
        RECT 95.215 79.175 95.505 79.345 ;
        RECT 95.675 79.175 95.965 79.345 ;
        RECT 96.135 79.175 96.425 79.345 ;
        RECT 96.595 79.175 96.885 79.345 ;
        RECT 97.055 79.175 97.345 79.345 ;
        RECT 97.515 79.175 97.805 79.345 ;
        RECT 97.975 79.175 98.265 79.345 ;
        RECT 98.435 79.175 98.725 79.345 ;
        RECT 98.895 79.175 99.185 79.345 ;
        RECT 99.355 79.175 99.645 79.345 ;
        RECT 99.815 79.175 99.960 79.345 ;
        RECT 16.785 78.425 17.995 79.175 ;
        RECT 16.785 77.885 17.305 78.425 ;
        RECT 18.165 78.405 23.510 79.175 ;
        RECT 23.685 78.405 29.030 79.175 ;
        RECT 29.205 78.405 30.875 79.175 ;
        RECT 31.045 78.450 31.335 79.175 ;
        RECT 31.505 78.405 36.850 79.175 ;
        RECT 37.025 78.405 38.695 79.175 ;
        RECT 38.955 78.625 39.125 78.915 ;
        RECT 39.295 78.795 39.625 79.175 ;
        RECT 38.955 78.455 39.620 78.625 ;
        RECT 17.475 77.715 17.995 78.255 ;
        RECT 18.165 77.885 20.745 78.405 ;
        RECT 20.915 77.715 23.510 78.235 ;
        RECT 23.685 77.885 26.265 78.405 ;
        RECT 26.435 77.715 29.030 78.235 ;
        RECT 29.205 77.885 29.955 78.405 ;
        RECT 30.125 77.715 30.875 78.235 ;
        RECT 31.505 77.885 34.085 78.405 ;
        RECT 16.785 76.625 17.995 77.715 ;
        RECT 18.165 76.625 23.510 77.715 ;
        RECT 23.685 76.625 29.030 77.715 ;
        RECT 29.205 76.625 30.875 77.715 ;
        RECT 31.045 76.625 31.335 77.790 ;
        RECT 34.255 77.715 36.850 78.235 ;
        RECT 37.025 77.885 37.775 78.405 ;
        RECT 37.945 77.715 38.695 78.235 ;
        RECT 31.505 76.625 36.850 77.715 ;
        RECT 37.025 76.625 38.695 77.715 ;
      LAYER li1 ;
        RECT 38.870 77.635 39.220 78.285 ;
      LAYER li1 ;
        RECT 39.390 77.465 39.620 78.455 ;
        RECT 38.955 77.295 39.620 77.465 ;
        RECT 38.955 76.795 39.125 77.295 ;
        RECT 39.295 76.625 39.625 77.125 ;
        RECT 39.795 76.795 40.020 78.915 ;
        RECT 40.235 78.715 40.485 79.175 ;
        RECT 40.670 78.725 41.000 78.895 ;
        RECT 41.180 78.725 41.930 78.895 ;
      LAYER li1 ;
        RECT 40.220 77.595 40.500 78.195 ;
      LAYER li1 ;
        RECT 40.670 77.195 40.840 78.725 ;
        RECT 41.010 78.225 41.590 78.555 ;
        RECT 41.010 77.355 41.250 78.225 ;
        RECT 41.760 77.945 41.930 78.725 ;
        RECT 42.180 78.675 42.550 79.175 ;
        RECT 42.730 78.725 43.190 78.895 ;
        RECT 43.420 78.725 44.090 78.895 ;
        RECT 42.730 78.495 42.900 78.725 ;
        RECT 42.100 78.195 42.900 78.495 ;
        RECT 43.070 78.225 43.620 78.555 ;
        RECT 42.100 78.165 42.270 78.195 ;
        RECT 42.390 77.945 42.560 78.015 ;
        RECT 41.760 77.775 42.560 77.945 ;
        RECT 42.050 77.685 42.560 77.775 ;
        RECT 41.440 77.250 41.880 77.605 ;
        RECT 40.220 76.625 40.485 77.085 ;
        RECT 40.670 76.820 40.905 77.195 ;
        RECT 42.050 77.070 42.220 77.685 ;
        RECT 41.150 76.900 42.220 77.070 ;
        RECT 42.390 76.625 42.560 77.425 ;
        RECT 42.730 77.125 42.900 78.195 ;
        RECT 43.070 77.295 43.260 78.015 ;
        RECT 43.430 77.685 43.620 78.225 ;
        RECT 43.920 78.185 44.090 78.725 ;
        RECT 44.405 78.645 44.575 79.175 ;
        RECT 44.870 78.525 45.230 78.965 ;
        RECT 45.405 78.695 45.575 79.175 ;
        RECT 46.275 78.700 46.445 79.175 ;
        RECT 47.125 78.700 47.295 79.175 ;
        RECT 44.870 78.355 45.370 78.525 ;
        RECT 45.200 78.185 45.370 78.355 ;
        RECT 47.605 78.405 52.950 79.175 ;
        RECT 53.125 78.405 58.470 79.175 ;
        RECT 59.105 78.450 59.395 79.175 ;
        RECT 59.565 78.405 64.910 79.175 ;
        RECT 65.085 78.405 70.430 79.175 ;
        RECT 70.605 78.405 73.195 79.175 ;
        RECT 73.455 78.625 73.625 78.915 ;
        RECT 73.795 78.795 74.125 79.175 ;
        RECT 73.455 78.455 74.120 78.625 ;
        RECT 43.920 78.015 45.010 78.185 ;
        RECT 45.200 78.015 47.020 78.185 ;
        RECT 43.430 77.355 43.750 77.685 ;
        RECT 42.730 76.795 42.980 77.125 ;
        RECT 43.920 77.095 44.090 78.015 ;
        RECT 45.200 77.760 45.370 78.015 ;
        RECT 47.605 77.885 50.185 78.405 ;
        RECT 44.260 77.590 45.370 77.760 ;
        RECT 50.355 77.715 52.950 78.235 ;
        RECT 53.125 77.885 55.705 78.405 ;
        RECT 55.875 77.715 58.470 78.235 ;
        RECT 59.565 77.885 62.145 78.405 ;
        RECT 44.260 77.430 45.120 77.590 ;
        RECT 43.205 76.925 44.090 77.095 ;
        RECT 44.270 76.625 44.485 77.125 ;
        RECT 44.950 76.805 45.120 77.430 ;
        RECT 45.405 76.625 45.585 77.405 ;
        RECT 46.280 76.625 46.450 77.455 ;
        RECT 47.120 76.625 47.290 77.455 ;
        RECT 47.605 76.625 52.950 77.715 ;
        RECT 53.125 76.625 58.470 77.715 ;
        RECT 59.105 76.625 59.395 77.790 ;
        RECT 62.315 77.715 64.910 78.235 ;
        RECT 65.085 77.885 67.665 78.405 ;
        RECT 67.835 77.715 70.430 78.235 ;
        RECT 70.605 77.885 71.815 78.405 ;
        RECT 71.985 77.715 73.195 78.235 ;
        RECT 59.565 76.625 64.910 77.715 ;
        RECT 65.085 76.625 70.430 77.715 ;
        RECT 70.605 76.625 73.195 77.715 ;
      LAYER li1 ;
        RECT 73.370 77.635 73.720 78.285 ;
      LAYER li1 ;
        RECT 73.890 77.465 74.120 78.455 ;
        RECT 73.455 77.295 74.120 77.465 ;
        RECT 73.455 76.795 73.625 77.295 ;
        RECT 73.795 76.625 74.125 77.125 ;
        RECT 74.295 76.795 74.520 78.915 ;
        RECT 74.735 78.715 74.985 79.175 ;
        RECT 75.170 78.725 75.500 78.895 ;
        RECT 75.680 78.725 76.430 78.895 ;
      LAYER li1 ;
        RECT 74.720 77.595 75.000 78.195 ;
      LAYER li1 ;
        RECT 75.170 77.195 75.340 78.725 ;
        RECT 75.510 78.225 76.090 78.555 ;
        RECT 75.510 77.355 75.750 78.225 ;
        RECT 76.260 77.945 76.430 78.725 ;
        RECT 76.680 78.675 77.050 79.175 ;
        RECT 77.230 78.725 77.690 78.895 ;
        RECT 77.920 78.725 78.590 78.895 ;
        RECT 77.230 78.495 77.400 78.725 ;
        RECT 76.600 78.195 77.400 78.495 ;
        RECT 77.570 78.225 78.120 78.555 ;
        RECT 76.600 78.165 76.770 78.195 ;
        RECT 76.890 77.945 77.060 78.015 ;
        RECT 76.260 77.775 77.060 77.945 ;
        RECT 76.550 77.685 77.060 77.775 ;
        RECT 75.940 77.250 76.380 77.605 ;
        RECT 74.720 76.625 74.985 77.085 ;
        RECT 75.170 76.820 75.405 77.195 ;
        RECT 76.550 77.070 76.720 77.685 ;
        RECT 75.650 76.900 76.720 77.070 ;
        RECT 76.890 76.625 77.060 77.425 ;
        RECT 77.230 77.125 77.400 78.195 ;
        RECT 77.570 77.295 77.760 78.015 ;
        RECT 77.930 77.685 78.120 78.225 ;
        RECT 78.420 78.185 78.590 78.725 ;
        RECT 78.905 78.645 79.075 79.175 ;
        RECT 79.370 78.525 79.730 78.965 ;
        RECT 79.905 78.695 80.075 79.175 ;
        RECT 80.775 78.700 80.945 79.175 ;
        RECT 81.625 78.700 81.795 79.175 ;
        RECT 79.370 78.355 79.870 78.525 ;
        RECT 79.700 78.185 79.870 78.355 ;
        RECT 82.105 78.405 85.615 79.175 ;
        RECT 85.785 78.425 86.995 79.175 ;
        RECT 87.165 78.450 87.455 79.175 ;
        RECT 78.420 78.015 79.510 78.185 ;
        RECT 79.700 78.015 81.520 78.185 ;
        RECT 77.930 77.355 78.250 77.685 ;
        RECT 77.230 76.795 77.480 77.125 ;
        RECT 78.420 77.095 78.590 78.015 ;
        RECT 79.700 77.760 79.870 78.015 ;
        RECT 82.105 77.885 83.755 78.405 ;
        RECT 78.760 77.590 79.870 77.760 ;
        RECT 83.925 77.715 85.615 78.235 ;
        RECT 85.785 77.885 86.305 78.425 ;
        RECT 87.625 78.405 92.970 79.175 ;
        RECT 93.145 78.405 98.490 79.175 ;
        RECT 98.665 78.425 99.875 79.175 ;
        RECT 86.475 77.715 86.995 78.255 ;
        RECT 87.625 77.885 90.205 78.405 ;
        RECT 78.760 77.430 79.620 77.590 ;
        RECT 77.705 76.925 78.590 77.095 ;
        RECT 78.770 76.625 78.985 77.125 ;
        RECT 79.450 76.805 79.620 77.430 ;
        RECT 79.905 76.625 80.085 77.405 ;
        RECT 80.780 76.625 80.950 77.455 ;
        RECT 81.620 76.625 81.790 77.455 ;
        RECT 82.105 76.625 85.615 77.715 ;
        RECT 85.785 76.625 86.995 77.715 ;
        RECT 87.165 76.625 87.455 77.790 ;
        RECT 90.375 77.715 92.970 78.235 ;
        RECT 93.145 77.885 95.725 78.405 ;
        RECT 95.895 77.715 98.490 78.235 ;
        RECT 87.625 76.625 92.970 77.715 ;
        RECT 93.145 76.625 98.490 77.715 ;
        RECT 98.665 77.715 99.185 78.255 ;
        RECT 99.355 77.885 99.875 78.425 ;
        RECT 98.665 76.625 99.875 77.715 ;
        RECT 16.700 76.455 16.845 76.625 ;
        RECT 17.015 76.455 17.305 76.625 ;
        RECT 17.475 76.455 17.765 76.625 ;
        RECT 17.935 76.455 18.225 76.625 ;
        RECT 18.395 76.455 18.685 76.625 ;
        RECT 18.855 76.455 19.145 76.625 ;
        RECT 19.315 76.455 19.605 76.625 ;
        RECT 19.775 76.455 20.065 76.625 ;
        RECT 20.235 76.455 20.525 76.625 ;
        RECT 20.695 76.455 20.985 76.625 ;
        RECT 21.155 76.455 21.445 76.625 ;
        RECT 21.615 76.455 21.905 76.625 ;
        RECT 22.075 76.455 22.365 76.625 ;
        RECT 22.535 76.455 22.825 76.625 ;
        RECT 22.995 76.455 23.285 76.625 ;
        RECT 23.455 76.455 23.745 76.625 ;
        RECT 23.915 76.455 24.205 76.625 ;
        RECT 24.375 76.455 24.665 76.625 ;
        RECT 24.835 76.455 25.125 76.625 ;
        RECT 25.295 76.455 25.585 76.625 ;
        RECT 25.755 76.455 26.045 76.625 ;
        RECT 26.215 76.455 26.505 76.625 ;
        RECT 26.675 76.455 26.965 76.625 ;
        RECT 27.135 76.455 27.425 76.625 ;
        RECT 27.595 76.455 27.885 76.625 ;
        RECT 28.055 76.455 28.345 76.625 ;
        RECT 28.515 76.455 28.805 76.625 ;
        RECT 28.975 76.455 29.265 76.625 ;
        RECT 29.435 76.455 29.725 76.625 ;
        RECT 29.895 76.455 30.185 76.625 ;
        RECT 30.355 76.455 30.645 76.625 ;
        RECT 30.815 76.455 31.105 76.625 ;
        RECT 31.275 76.455 31.565 76.625 ;
        RECT 31.735 76.455 32.025 76.625 ;
        RECT 32.195 76.455 32.485 76.625 ;
        RECT 32.655 76.455 32.945 76.625 ;
        RECT 33.115 76.455 33.405 76.625 ;
        RECT 33.575 76.455 33.865 76.625 ;
        RECT 34.035 76.455 34.325 76.625 ;
        RECT 34.495 76.455 34.785 76.625 ;
        RECT 34.955 76.455 35.245 76.625 ;
        RECT 35.415 76.455 35.705 76.625 ;
        RECT 35.875 76.455 36.165 76.625 ;
        RECT 36.335 76.455 36.625 76.625 ;
        RECT 36.795 76.455 37.085 76.625 ;
        RECT 37.255 76.455 37.545 76.625 ;
        RECT 37.715 76.455 38.005 76.625 ;
        RECT 38.175 76.455 38.465 76.625 ;
        RECT 38.635 76.455 38.925 76.625 ;
        RECT 39.095 76.455 39.385 76.625 ;
        RECT 39.555 76.455 39.845 76.625 ;
        RECT 40.015 76.455 40.305 76.625 ;
        RECT 40.475 76.455 40.765 76.625 ;
        RECT 40.935 76.455 41.225 76.625 ;
        RECT 41.395 76.455 41.685 76.625 ;
        RECT 41.855 76.455 42.145 76.625 ;
        RECT 42.315 76.455 42.605 76.625 ;
        RECT 42.775 76.455 43.065 76.625 ;
        RECT 43.235 76.455 43.525 76.625 ;
        RECT 43.695 76.455 43.985 76.625 ;
        RECT 44.155 76.455 44.445 76.625 ;
        RECT 44.615 76.455 44.905 76.625 ;
        RECT 45.075 76.455 45.365 76.625 ;
        RECT 45.535 76.455 45.825 76.625 ;
        RECT 45.995 76.455 46.285 76.625 ;
        RECT 46.455 76.455 46.745 76.625 ;
        RECT 46.915 76.455 47.205 76.625 ;
        RECT 47.375 76.455 47.665 76.625 ;
        RECT 47.835 76.455 48.125 76.625 ;
        RECT 48.295 76.455 48.585 76.625 ;
        RECT 48.755 76.455 49.045 76.625 ;
        RECT 49.215 76.455 49.505 76.625 ;
        RECT 49.675 76.455 49.965 76.625 ;
        RECT 50.135 76.455 50.425 76.625 ;
        RECT 50.595 76.455 50.885 76.625 ;
        RECT 51.055 76.455 51.345 76.625 ;
        RECT 51.515 76.455 51.805 76.625 ;
        RECT 51.975 76.455 52.265 76.625 ;
        RECT 52.435 76.455 52.725 76.625 ;
        RECT 52.895 76.455 53.185 76.625 ;
        RECT 53.355 76.455 53.645 76.625 ;
        RECT 53.815 76.455 54.105 76.625 ;
        RECT 54.275 76.455 54.565 76.625 ;
        RECT 54.735 76.455 55.025 76.625 ;
        RECT 55.195 76.455 55.485 76.625 ;
        RECT 55.655 76.455 55.945 76.625 ;
        RECT 56.115 76.455 56.405 76.625 ;
        RECT 56.575 76.455 56.865 76.625 ;
        RECT 57.035 76.455 57.325 76.625 ;
        RECT 57.495 76.455 57.785 76.625 ;
        RECT 57.955 76.455 58.245 76.625 ;
        RECT 58.415 76.455 58.705 76.625 ;
        RECT 58.875 76.455 59.165 76.625 ;
        RECT 59.335 76.455 59.625 76.625 ;
        RECT 59.795 76.455 60.085 76.625 ;
        RECT 60.255 76.455 60.545 76.625 ;
        RECT 60.715 76.455 61.005 76.625 ;
        RECT 61.175 76.455 61.465 76.625 ;
        RECT 61.635 76.455 61.925 76.625 ;
        RECT 62.095 76.455 62.385 76.625 ;
        RECT 62.555 76.455 62.845 76.625 ;
        RECT 63.015 76.455 63.305 76.625 ;
        RECT 63.475 76.455 63.765 76.625 ;
        RECT 63.935 76.455 64.225 76.625 ;
        RECT 64.395 76.455 64.685 76.625 ;
        RECT 64.855 76.455 65.145 76.625 ;
        RECT 65.315 76.455 65.605 76.625 ;
        RECT 65.775 76.455 66.065 76.625 ;
        RECT 66.235 76.455 66.525 76.625 ;
        RECT 66.695 76.455 66.985 76.625 ;
        RECT 67.155 76.455 67.445 76.625 ;
        RECT 67.615 76.455 67.905 76.625 ;
        RECT 68.075 76.455 68.365 76.625 ;
        RECT 68.535 76.455 68.825 76.625 ;
        RECT 68.995 76.455 69.285 76.625 ;
        RECT 69.455 76.455 69.745 76.625 ;
        RECT 69.915 76.455 70.205 76.625 ;
        RECT 70.375 76.455 70.665 76.625 ;
        RECT 70.835 76.455 71.125 76.625 ;
        RECT 71.295 76.455 71.585 76.625 ;
        RECT 71.755 76.455 72.045 76.625 ;
        RECT 72.215 76.455 72.505 76.625 ;
        RECT 72.675 76.455 72.965 76.625 ;
        RECT 73.135 76.455 73.425 76.625 ;
        RECT 73.595 76.455 73.885 76.625 ;
        RECT 74.055 76.455 74.345 76.625 ;
        RECT 74.515 76.455 74.805 76.625 ;
        RECT 74.975 76.455 75.265 76.625 ;
        RECT 75.435 76.455 75.725 76.625 ;
        RECT 75.895 76.455 76.185 76.625 ;
        RECT 76.355 76.455 76.645 76.625 ;
        RECT 76.815 76.455 77.105 76.625 ;
        RECT 77.275 76.455 77.565 76.625 ;
        RECT 77.735 76.455 78.025 76.625 ;
        RECT 78.195 76.455 78.485 76.625 ;
        RECT 78.655 76.455 78.945 76.625 ;
        RECT 79.115 76.455 79.405 76.625 ;
        RECT 79.575 76.455 79.865 76.625 ;
        RECT 80.035 76.455 80.325 76.625 ;
        RECT 80.495 76.455 80.785 76.625 ;
        RECT 80.955 76.455 81.245 76.625 ;
        RECT 81.415 76.455 81.705 76.625 ;
        RECT 81.875 76.455 82.165 76.625 ;
        RECT 82.335 76.455 82.625 76.625 ;
        RECT 82.795 76.455 83.085 76.625 ;
        RECT 83.255 76.455 83.545 76.625 ;
        RECT 83.715 76.455 84.005 76.625 ;
        RECT 84.175 76.455 84.465 76.625 ;
        RECT 84.635 76.455 84.925 76.625 ;
        RECT 85.095 76.455 85.385 76.625 ;
        RECT 85.555 76.455 85.845 76.625 ;
        RECT 86.015 76.455 86.305 76.625 ;
        RECT 86.475 76.455 86.765 76.625 ;
        RECT 86.935 76.455 87.225 76.625 ;
        RECT 87.395 76.455 87.685 76.625 ;
        RECT 87.855 76.455 88.145 76.625 ;
        RECT 88.315 76.455 88.605 76.625 ;
        RECT 88.775 76.455 89.065 76.625 ;
        RECT 89.235 76.455 89.525 76.625 ;
        RECT 89.695 76.455 89.985 76.625 ;
        RECT 90.155 76.455 90.445 76.625 ;
        RECT 90.615 76.455 90.905 76.625 ;
        RECT 91.075 76.455 91.365 76.625 ;
        RECT 91.535 76.455 91.825 76.625 ;
        RECT 91.995 76.455 92.285 76.625 ;
        RECT 92.455 76.455 92.745 76.625 ;
        RECT 92.915 76.455 93.205 76.625 ;
        RECT 93.375 76.455 93.665 76.625 ;
        RECT 93.835 76.455 94.125 76.625 ;
        RECT 94.295 76.455 94.585 76.625 ;
        RECT 94.755 76.455 95.045 76.625 ;
        RECT 95.215 76.455 95.505 76.625 ;
        RECT 95.675 76.455 95.965 76.625 ;
        RECT 96.135 76.455 96.425 76.625 ;
        RECT 96.595 76.455 96.885 76.625 ;
        RECT 97.055 76.455 97.345 76.625 ;
        RECT 97.515 76.455 97.805 76.625 ;
        RECT 97.975 76.455 98.265 76.625 ;
        RECT 98.435 76.455 98.725 76.625 ;
        RECT 98.895 76.455 99.185 76.625 ;
        RECT 99.355 76.455 99.645 76.625 ;
        RECT 99.815 76.455 99.960 76.625 ;
        RECT 16.785 75.365 17.995 76.455 ;
        RECT 18.165 75.365 23.510 76.455 ;
        RECT 23.685 75.365 29.030 76.455 ;
        RECT 29.205 75.365 34.550 76.455 ;
        RECT 34.725 75.365 40.070 76.455 ;
        RECT 40.245 75.365 43.755 76.455 ;
        RECT 16.785 74.655 17.305 75.195 ;
        RECT 17.475 74.825 17.995 75.365 ;
        RECT 18.165 74.675 20.745 75.195 ;
        RECT 20.915 74.845 23.510 75.365 ;
        RECT 23.685 74.675 26.265 75.195 ;
        RECT 26.435 74.845 29.030 75.365 ;
        RECT 29.205 74.675 31.785 75.195 ;
        RECT 31.955 74.845 34.550 75.365 ;
        RECT 34.725 74.675 37.305 75.195 ;
        RECT 37.475 74.845 40.070 75.365 ;
        RECT 40.245 74.675 41.895 75.195 ;
        RECT 42.065 74.845 43.755 75.365 ;
        RECT 44.845 75.290 45.135 76.455 ;
        RECT 45.305 75.365 50.650 76.455 ;
        RECT 50.825 75.365 56.170 76.455 ;
        RECT 56.345 75.365 61.690 76.455 ;
        RECT 61.865 75.365 67.210 76.455 ;
        RECT 67.385 75.365 72.730 76.455 ;
        RECT 45.305 74.675 47.885 75.195 ;
        RECT 48.055 74.845 50.650 75.365 ;
        RECT 50.825 74.675 53.405 75.195 ;
        RECT 53.575 74.845 56.170 75.365 ;
        RECT 56.345 74.675 58.925 75.195 ;
        RECT 59.095 74.845 61.690 75.365 ;
        RECT 61.865 74.675 64.445 75.195 ;
        RECT 64.615 74.845 67.210 75.365 ;
        RECT 67.385 74.675 69.965 75.195 ;
        RECT 70.135 74.845 72.730 75.365 ;
        RECT 72.905 75.290 73.195 76.455 ;
        RECT 73.365 75.365 78.710 76.455 ;
        RECT 78.885 75.365 84.230 76.455 ;
        RECT 84.405 75.365 89.750 76.455 ;
        RECT 89.925 75.365 95.270 76.455 ;
        RECT 95.445 75.365 98.035 76.455 ;
        RECT 73.365 74.675 75.945 75.195 ;
        RECT 76.115 74.845 78.710 75.365 ;
        RECT 78.885 74.675 81.465 75.195 ;
        RECT 81.635 74.845 84.230 75.365 ;
        RECT 84.405 74.675 86.985 75.195 ;
        RECT 87.155 74.845 89.750 75.365 ;
        RECT 89.925 74.675 92.505 75.195 ;
        RECT 92.675 74.845 95.270 75.365 ;
        RECT 95.445 74.675 96.655 75.195 ;
        RECT 96.825 74.845 98.035 75.365 ;
        RECT 98.665 75.365 99.875 76.455 ;
        RECT 98.665 74.825 99.185 75.365 ;
        RECT 16.785 73.905 17.995 74.655 ;
        RECT 18.165 73.905 23.510 74.675 ;
        RECT 23.685 73.905 29.030 74.675 ;
        RECT 29.205 73.905 34.550 74.675 ;
        RECT 34.725 73.905 40.070 74.675 ;
        RECT 40.245 73.905 43.755 74.675 ;
        RECT 44.845 73.905 45.135 74.630 ;
        RECT 45.305 73.905 50.650 74.675 ;
        RECT 50.825 73.905 56.170 74.675 ;
        RECT 56.345 73.905 61.690 74.675 ;
        RECT 61.865 73.905 67.210 74.675 ;
        RECT 67.385 73.905 72.730 74.675 ;
        RECT 72.905 73.905 73.195 74.630 ;
        RECT 73.365 73.905 78.710 74.675 ;
        RECT 78.885 73.905 84.230 74.675 ;
        RECT 84.405 73.905 89.750 74.675 ;
        RECT 89.925 73.905 95.270 74.675 ;
        RECT 95.445 73.905 98.035 74.675 ;
        RECT 99.355 74.655 99.875 75.195 ;
        RECT 98.665 73.905 99.875 74.655 ;
        RECT 16.700 73.735 16.845 73.905 ;
        RECT 17.015 73.735 17.305 73.905 ;
        RECT 17.475 73.735 17.765 73.905 ;
        RECT 17.935 73.735 18.225 73.905 ;
        RECT 18.395 73.735 18.685 73.905 ;
        RECT 18.855 73.735 19.145 73.905 ;
        RECT 19.315 73.735 19.605 73.905 ;
        RECT 19.775 73.735 20.065 73.905 ;
        RECT 20.235 73.735 20.525 73.905 ;
        RECT 20.695 73.735 20.985 73.905 ;
        RECT 21.155 73.735 21.445 73.905 ;
        RECT 21.615 73.735 21.905 73.905 ;
        RECT 22.075 73.735 22.365 73.905 ;
        RECT 22.535 73.735 22.825 73.905 ;
        RECT 22.995 73.735 23.285 73.905 ;
        RECT 23.455 73.735 23.745 73.905 ;
        RECT 23.915 73.735 24.205 73.905 ;
        RECT 24.375 73.735 24.665 73.905 ;
        RECT 24.835 73.735 25.125 73.905 ;
        RECT 25.295 73.735 25.585 73.905 ;
        RECT 25.755 73.735 26.045 73.905 ;
        RECT 26.215 73.735 26.505 73.905 ;
        RECT 26.675 73.735 26.965 73.905 ;
        RECT 27.135 73.735 27.425 73.905 ;
        RECT 27.595 73.735 27.885 73.905 ;
        RECT 28.055 73.735 28.345 73.905 ;
        RECT 28.515 73.735 28.805 73.905 ;
        RECT 28.975 73.735 29.265 73.905 ;
        RECT 29.435 73.735 29.725 73.905 ;
        RECT 29.895 73.735 30.185 73.905 ;
        RECT 30.355 73.735 30.645 73.905 ;
        RECT 30.815 73.735 31.105 73.905 ;
        RECT 31.275 73.735 31.565 73.905 ;
        RECT 31.735 73.735 32.025 73.905 ;
        RECT 32.195 73.735 32.485 73.905 ;
        RECT 32.655 73.735 32.945 73.905 ;
        RECT 33.115 73.735 33.405 73.905 ;
        RECT 33.575 73.735 33.865 73.905 ;
        RECT 34.035 73.735 34.325 73.905 ;
        RECT 34.495 73.735 34.785 73.905 ;
        RECT 34.955 73.735 35.245 73.905 ;
        RECT 35.415 73.735 35.705 73.905 ;
        RECT 35.875 73.735 36.165 73.905 ;
        RECT 36.335 73.735 36.625 73.905 ;
        RECT 36.795 73.735 37.085 73.905 ;
        RECT 37.255 73.735 37.545 73.905 ;
        RECT 37.715 73.735 38.005 73.905 ;
        RECT 38.175 73.735 38.465 73.905 ;
        RECT 38.635 73.735 38.925 73.905 ;
        RECT 39.095 73.735 39.385 73.905 ;
        RECT 39.555 73.735 39.845 73.905 ;
        RECT 40.015 73.735 40.305 73.905 ;
        RECT 40.475 73.735 40.765 73.905 ;
        RECT 40.935 73.735 41.225 73.905 ;
        RECT 41.395 73.735 41.685 73.905 ;
        RECT 41.855 73.735 42.145 73.905 ;
        RECT 42.315 73.735 42.605 73.905 ;
        RECT 42.775 73.735 43.065 73.905 ;
        RECT 43.235 73.735 43.525 73.905 ;
        RECT 43.695 73.735 43.985 73.905 ;
        RECT 44.155 73.735 44.445 73.905 ;
        RECT 44.615 73.735 44.905 73.905 ;
        RECT 45.075 73.735 45.365 73.905 ;
        RECT 45.535 73.735 45.825 73.905 ;
        RECT 45.995 73.735 46.285 73.905 ;
        RECT 46.455 73.735 46.745 73.905 ;
        RECT 46.915 73.735 47.205 73.905 ;
        RECT 47.375 73.735 47.665 73.905 ;
        RECT 47.835 73.735 48.125 73.905 ;
        RECT 48.295 73.735 48.585 73.905 ;
        RECT 48.755 73.735 49.045 73.905 ;
        RECT 49.215 73.735 49.505 73.905 ;
        RECT 49.675 73.735 49.965 73.905 ;
        RECT 50.135 73.735 50.425 73.905 ;
        RECT 50.595 73.735 50.885 73.905 ;
        RECT 51.055 73.735 51.345 73.905 ;
        RECT 51.515 73.735 51.805 73.905 ;
        RECT 51.975 73.735 52.265 73.905 ;
        RECT 52.435 73.735 52.725 73.905 ;
        RECT 52.895 73.735 53.185 73.905 ;
        RECT 53.355 73.735 53.645 73.905 ;
        RECT 53.815 73.735 54.105 73.905 ;
        RECT 54.275 73.735 54.565 73.905 ;
        RECT 54.735 73.735 55.025 73.905 ;
        RECT 55.195 73.735 55.485 73.905 ;
        RECT 55.655 73.735 55.945 73.905 ;
        RECT 56.115 73.735 56.405 73.905 ;
        RECT 56.575 73.735 56.865 73.905 ;
        RECT 57.035 73.735 57.325 73.905 ;
        RECT 57.495 73.735 57.785 73.905 ;
        RECT 57.955 73.735 58.245 73.905 ;
        RECT 58.415 73.735 58.705 73.905 ;
        RECT 58.875 73.735 59.165 73.905 ;
        RECT 59.335 73.735 59.625 73.905 ;
        RECT 59.795 73.735 60.085 73.905 ;
        RECT 60.255 73.735 60.545 73.905 ;
        RECT 60.715 73.735 61.005 73.905 ;
        RECT 61.175 73.735 61.465 73.905 ;
        RECT 61.635 73.735 61.925 73.905 ;
        RECT 62.095 73.735 62.385 73.905 ;
        RECT 62.555 73.735 62.845 73.905 ;
        RECT 63.015 73.735 63.305 73.905 ;
        RECT 63.475 73.735 63.765 73.905 ;
        RECT 63.935 73.735 64.225 73.905 ;
        RECT 64.395 73.735 64.685 73.905 ;
        RECT 64.855 73.735 65.145 73.905 ;
        RECT 65.315 73.735 65.605 73.905 ;
        RECT 65.775 73.735 66.065 73.905 ;
        RECT 66.235 73.735 66.525 73.905 ;
        RECT 66.695 73.735 66.985 73.905 ;
        RECT 67.155 73.735 67.445 73.905 ;
        RECT 67.615 73.735 67.905 73.905 ;
        RECT 68.075 73.735 68.365 73.905 ;
        RECT 68.535 73.735 68.825 73.905 ;
        RECT 68.995 73.735 69.285 73.905 ;
        RECT 69.455 73.735 69.745 73.905 ;
        RECT 69.915 73.735 70.205 73.905 ;
        RECT 70.375 73.735 70.665 73.905 ;
        RECT 70.835 73.735 71.125 73.905 ;
        RECT 71.295 73.735 71.585 73.905 ;
        RECT 71.755 73.735 72.045 73.905 ;
        RECT 72.215 73.735 72.505 73.905 ;
        RECT 72.675 73.735 72.965 73.905 ;
        RECT 73.135 73.735 73.425 73.905 ;
        RECT 73.595 73.735 73.885 73.905 ;
        RECT 74.055 73.735 74.345 73.905 ;
        RECT 74.515 73.735 74.805 73.905 ;
        RECT 74.975 73.735 75.265 73.905 ;
        RECT 75.435 73.735 75.725 73.905 ;
        RECT 75.895 73.735 76.185 73.905 ;
        RECT 76.355 73.735 76.645 73.905 ;
        RECT 76.815 73.735 77.105 73.905 ;
        RECT 77.275 73.735 77.565 73.905 ;
        RECT 77.735 73.735 78.025 73.905 ;
        RECT 78.195 73.735 78.485 73.905 ;
        RECT 78.655 73.735 78.945 73.905 ;
        RECT 79.115 73.735 79.405 73.905 ;
        RECT 79.575 73.735 79.865 73.905 ;
        RECT 80.035 73.735 80.325 73.905 ;
        RECT 80.495 73.735 80.785 73.905 ;
        RECT 80.955 73.735 81.245 73.905 ;
        RECT 81.415 73.735 81.705 73.905 ;
        RECT 81.875 73.735 82.165 73.905 ;
        RECT 82.335 73.735 82.625 73.905 ;
        RECT 82.795 73.735 83.085 73.905 ;
        RECT 83.255 73.735 83.545 73.905 ;
        RECT 83.715 73.735 84.005 73.905 ;
        RECT 84.175 73.735 84.465 73.905 ;
        RECT 84.635 73.735 84.925 73.905 ;
        RECT 85.095 73.735 85.385 73.905 ;
        RECT 85.555 73.735 85.845 73.905 ;
        RECT 86.015 73.735 86.305 73.905 ;
        RECT 86.475 73.735 86.765 73.905 ;
        RECT 86.935 73.735 87.225 73.905 ;
        RECT 87.395 73.735 87.685 73.905 ;
        RECT 87.855 73.735 88.145 73.905 ;
        RECT 88.315 73.735 88.605 73.905 ;
        RECT 88.775 73.735 89.065 73.905 ;
        RECT 89.235 73.735 89.525 73.905 ;
        RECT 89.695 73.735 89.985 73.905 ;
        RECT 90.155 73.735 90.445 73.905 ;
        RECT 90.615 73.735 90.905 73.905 ;
        RECT 91.075 73.735 91.365 73.905 ;
        RECT 91.535 73.735 91.825 73.905 ;
        RECT 91.995 73.735 92.285 73.905 ;
        RECT 92.455 73.735 92.745 73.905 ;
        RECT 92.915 73.735 93.205 73.905 ;
        RECT 93.375 73.735 93.665 73.905 ;
        RECT 93.835 73.735 94.125 73.905 ;
        RECT 94.295 73.735 94.585 73.905 ;
        RECT 94.755 73.735 95.045 73.905 ;
        RECT 95.215 73.735 95.505 73.905 ;
        RECT 95.675 73.735 95.965 73.905 ;
        RECT 96.135 73.735 96.425 73.905 ;
        RECT 96.595 73.735 96.885 73.905 ;
        RECT 97.055 73.735 97.345 73.905 ;
        RECT 97.515 73.735 97.805 73.905 ;
        RECT 97.975 73.735 98.265 73.905 ;
        RECT 98.435 73.735 98.725 73.905 ;
        RECT 98.895 73.735 99.185 73.905 ;
        RECT 99.355 73.735 99.645 73.905 ;
        RECT 99.815 73.735 99.960 73.905 ;
        RECT 16.785 72.985 17.995 73.735 ;
        RECT 16.785 72.445 17.305 72.985 ;
        RECT 18.165 72.965 23.510 73.735 ;
        RECT 23.685 72.965 29.030 73.735 ;
        RECT 29.205 72.965 30.875 73.735 ;
        RECT 31.045 73.010 31.335 73.735 ;
        RECT 31.505 72.965 36.850 73.735 ;
        RECT 37.025 72.965 42.370 73.735 ;
        RECT 42.545 72.965 47.890 73.735 ;
        RECT 48.065 72.965 53.410 73.735 ;
        RECT 53.585 72.965 58.930 73.735 ;
        RECT 59.105 73.010 59.395 73.735 ;
        RECT 59.565 72.965 64.910 73.735 ;
        RECT 65.085 72.965 70.430 73.735 ;
        RECT 70.605 72.965 75.950 73.735 ;
        RECT 76.125 72.965 81.470 73.735 ;
        RECT 81.645 72.965 86.990 73.735 ;
        RECT 87.165 73.010 87.455 73.735 ;
        RECT 87.625 72.965 92.970 73.735 ;
        RECT 93.145 72.965 98.490 73.735 ;
        RECT 98.665 72.985 99.875 73.735 ;
        RECT 17.475 72.275 17.995 72.815 ;
        RECT 18.165 72.445 20.745 72.965 ;
        RECT 20.915 72.275 23.510 72.795 ;
        RECT 23.685 72.445 26.265 72.965 ;
        RECT 26.435 72.275 29.030 72.795 ;
        RECT 29.205 72.445 29.955 72.965 ;
        RECT 30.125 72.275 30.875 72.795 ;
        RECT 31.505 72.445 34.085 72.965 ;
        RECT 16.785 71.185 17.995 72.275 ;
        RECT 18.165 71.185 23.510 72.275 ;
        RECT 23.685 71.185 29.030 72.275 ;
        RECT 29.205 71.185 30.875 72.275 ;
        RECT 31.045 71.185 31.335 72.350 ;
        RECT 34.255 72.275 36.850 72.795 ;
        RECT 37.025 72.445 39.605 72.965 ;
        RECT 39.775 72.275 42.370 72.795 ;
        RECT 42.545 72.445 45.125 72.965 ;
        RECT 45.295 72.275 47.890 72.795 ;
        RECT 48.065 72.445 50.645 72.965 ;
        RECT 50.815 72.275 53.410 72.795 ;
        RECT 53.585 72.445 56.165 72.965 ;
        RECT 56.335 72.275 58.930 72.795 ;
        RECT 59.565 72.445 62.145 72.965 ;
        RECT 31.505 71.185 36.850 72.275 ;
        RECT 37.025 71.185 42.370 72.275 ;
        RECT 42.545 71.185 47.890 72.275 ;
        RECT 48.065 71.185 53.410 72.275 ;
        RECT 53.585 71.185 58.930 72.275 ;
        RECT 59.105 71.185 59.395 72.350 ;
        RECT 62.315 72.275 64.910 72.795 ;
        RECT 65.085 72.445 67.665 72.965 ;
        RECT 67.835 72.275 70.430 72.795 ;
        RECT 70.605 72.445 73.185 72.965 ;
        RECT 73.355 72.275 75.950 72.795 ;
        RECT 76.125 72.445 78.705 72.965 ;
        RECT 78.875 72.275 81.470 72.795 ;
        RECT 81.645 72.445 84.225 72.965 ;
        RECT 84.395 72.275 86.990 72.795 ;
        RECT 87.625 72.445 90.205 72.965 ;
        RECT 59.565 71.185 64.910 72.275 ;
        RECT 65.085 71.185 70.430 72.275 ;
        RECT 70.605 71.185 75.950 72.275 ;
        RECT 76.125 71.185 81.470 72.275 ;
        RECT 81.645 71.185 86.990 72.275 ;
        RECT 87.165 71.185 87.455 72.350 ;
        RECT 90.375 72.275 92.970 72.795 ;
        RECT 93.145 72.445 95.725 72.965 ;
        RECT 95.895 72.275 98.490 72.795 ;
        RECT 87.625 71.185 92.970 72.275 ;
        RECT 93.145 71.185 98.490 72.275 ;
        RECT 98.665 72.275 99.185 72.815 ;
        RECT 99.355 72.445 99.875 72.985 ;
        RECT 98.665 71.185 99.875 72.275 ;
        RECT 16.700 71.015 16.845 71.185 ;
        RECT 17.015 71.015 17.305 71.185 ;
        RECT 17.475 71.015 17.765 71.185 ;
        RECT 17.935 71.015 18.225 71.185 ;
        RECT 18.395 71.015 18.685 71.185 ;
        RECT 18.855 71.015 19.145 71.185 ;
        RECT 19.315 71.015 19.605 71.185 ;
        RECT 19.775 71.015 20.065 71.185 ;
        RECT 20.235 71.015 20.525 71.185 ;
        RECT 20.695 71.015 20.985 71.185 ;
        RECT 21.155 71.015 21.445 71.185 ;
        RECT 21.615 71.015 21.905 71.185 ;
        RECT 22.075 71.015 22.365 71.185 ;
        RECT 22.535 71.015 22.825 71.185 ;
        RECT 22.995 71.015 23.285 71.185 ;
        RECT 23.455 71.015 23.745 71.185 ;
        RECT 23.915 71.015 24.205 71.185 ;
        RECT 24.375 71.015 24.665 71.185 ;
        RECT 24.835 71.015 25.125 71.185 ;
        RECT 25.295 71.015 25.585 71.185 ;
        RECT 25.755 71.015 26.045 71.185 ;
        RECT 26.215 71.015 26.505 71.185 ;
        RECT 26.675 71.015 26.965 71.185 ;
        RECT 27.135 71.015 27.425 71.185 ;
        RECT 27.595 71.015 27.885 71.185 ;
        RECT 28.055 71.015 28.345 71.185 ;
        RECT 28.515 71.015 28.805 71.185 ;
        RECT 28.975 71.015 29.265 71.185 ;
        RECT 29.435 71.015 29.725 71.185 ;
        RECT 29.895 71.015 30.185 71.185 ;
        RECT 30.355 71.015 30.645 71.185 ;
        RECT 30.815 71.015 31.105 71.185 ;
        RECT 31.275 71.015 31.565 71.185 ;
        RECT 31.735 71.015 32.025 71.185 ;
        RECT 32.195 71.015 32.485 71.185 ;
        RECT 32.655 71.015 32.945 71.185 ;
        RECT 33.115 71.015 33.405 71.185 ;
        RECT 33.575 71.015 33.865 71.185 ;
        RECT 34.035 71.015 34.325 71.185 ;
        RECT 34.495 71.015 34.785 71.185 ;
        RECT 34.955 71.015 35.245 71.185 ;
        RECT 35.415 71.015 35.705 71.185 ;
        RECT 35.875 71.015 36.165 71.185 ;
        RECT 36.335 71.015 36.625 71.185 ;
        RECT 36.795 71.015 37.085 71.185 ;
        RECT 37.255 71.015 37.545 71.185 ;
        RECT 37.715 71.015 38.005 71.185 ;
        RECT 38.175 71.015 38.465 71.185 ;
        RECT 38.635 71.015 38.925 71.185 ;
        RECT 39.095 71.015 39.385 71.185 ;
        RECT 39.555 71.015 39.845 71.185 ;
        RECT 40.015 71.015 40.305 71.185 ;
        RECT 40.475 71.015 40.765 71.185 ;
        RECT 40.935 71.015 41.225 71.185 ;
        RECT 41.395 71.015 41.685 71.185 ;
        RECT 41.855 71.015 42.145 71.185 ;
        RECT 42.315 71.015 42.605 71.185 ;
        RECT 42.775 71.015 43.065 71.185 ;
        RECT 43.235 71.015 43.525 71.185 ;
        RECT 43.695 71.015 43.985 71.185 ;
        RECT 44.155 71.015 44.445 71.185 ;
        RECT 44.615 71.015 44.905 71.185 ;
        RECT 45.075 71.015 45.365 71.185 ;
        RECT 45.535 71.015 45.825 71.185 ;
        RECT 45.995 71.015 46.285 71.185 ;
        RECT 46.455 71.015 46.745 71.185 ;
        RECT 46.915 71.015 47.205 71.185 ;
        RECT 47.375 71.015 47.665 71.185 ;
        RECT 47.835 71.015 48.125 71.185 ;
        RECT 48.295 71.015 48.585 71.185 ;
        RECT 48.755 71.015 49.045 71.185 ;
        RECT 49.215 71.015 49.505 71.185 ;
        RECT 49.675 71.015 49.965 71.185 ;
        RECT 50.135 71.015 50.425 71.185 ;
        RECT 50.595 71.015 50.885 71.185 ;
        RECT 51.055 71.015 51.345 71.185 ;
        RECT 51.515 71.015 51.805 71.185 ;
        RECT 51.975 71.015 52.265 71.185 ;
        RECT 52.435 71.015 52.725 71.185 ;
        RECT 52.895 71.015 53.185 71.185 ;
        RECT 53.355 71.015 53.645 71.185 ;
        RECT 53.815 71.015 54.105 71.185 ;
        RECT 54.275 71.015 54.565 71.185 ;
        RECT 54.735 71.015 55.025 71.185 ;
        RECT 55.195 71.015 55.485 71.185 ;
        RECT 55.655 71.015 55.945 71.185 ;
        RECT 56.115 71.015 56.405 71.185 ;
        RECT 56.575 71.015 56.865 71.185 ;
        RECT 57.035 71.015 57.325 71.185 ;
        RECT 57.495 71.015 57.785 71.185 ;
        RECT 57.955 71.015 58.245 71.185 ;
        RECT 58.415 71.015 58.705 71.185 ;
        RECT 58.875 71.015 59.165 71.185 ;
        RECT 59.335 71.015 59.625 71.185 ;
        RECT 59.795 71.015 60.085 71.185 ;
        RECT 60.255 71.015 60.545 71.185 ;
        RECT 60.715 71.015 61.005 71.185 ;
        RECT 61.175 71.015 61.465 71.185 ;
        RECT 61.635 71.015 61.925 71.185 ;
        RECT 62.095 71.015 62.385 71.185 ;
        RECT 62.555 71.015 62.845 71.185 ;
        RECT 63.015 71.015 63.305 71.185 ;
        RECT 63.475 71.015 63.765 71.185 ;
        RECT 63.935 71.015 64.225 71.185 ;
        RECT 64.395 71.015 64.685 71.185 ;
        RECT 64.855 71.015 65.145 71.185 ;
        RECT 65.315 71.015 65.605 71.185 ;
        RECT 65.775 71.015 66.065 71.185 ;
        RECT 66.235 71.015 66.525 71.185 ;
        RECT 66.695 71.015 66.985 71.185 ;
        RECT 67.155 71.015 67.445 71.185 ;
        RECT 67.615 71.015 67.905 71.185 ;
        RECT 68.075 71.015 68.365 71.185 ;
        RECT 68.535 71.015 68.825 71.185 ;
        RECT 68.995 71.015 69.285 71.185 ;
        RECT 69.455 71.015 69.745 71.185 ;
        RECT 69.915 71.015 70.205 71.185 ;
        RECT 70.375 71.015 70.665 71.185 ;
        RECT 70.835 71.015 71.125 71.185 ;
        RECT 71.295 71.015 71.585 71.185 ;
        RECT 71.755 71.015 72.045 71.185 ;
        RECT 72.215 71.015 72.505 71.185 ;
        RECT 72.675 71.015 72.965 71.185 ;
        RECT 73.135 71.015 73.425 71.185 ;
        RECT 73.595 71.015 73.885 71.185 ;
        RECT 74.055 71.015 74.345 71.185 ;
        RECT 74.515 71.015 74.805 71.185 ;
        RECT 74.975 71.015 75.265 71.185 ;
        RECT 75.435 71.015 75.725 71.185 ;
        RECT 75.895 71.015 76.185 71.185 ;
        RECT 76.355 71.015 76.645 71.185 ;
        RECT 76.815 71.015 77.105 71.185 ;
        RECT 77.275 71.015 77.565 71.185 ;
        RECT 77.735 71.015 78.025 71.185 ;
        RECT 78.195 71.015 78.485 71.185 ;
        RECT 78.655 71.015 78.945 71.185 ;
        RECT 79.115 71.015 79.405 71.185 ;
        RECT 79.575 71.015 79.865 71.185 ;
        RECT 80.035 71.015 80.325 71.185 ;
        RECT 80.495 71.015 80.785 71.185 ;
        RECT 80.955 71.015 81.245 71.185 ;
        RECT 81.415 71.015 81.705 71.185 ;
        RECT 81.875 71.015 82.165 71.185 ;
        RECT 82.335 71.015 82.625 71.185 ;
        RECT 82.795 71.015 83.085 71.185 ;
        RECT 83.255 71.015 83.545 71.185 ;
        RECT 83.715 71.015 84.005 71.185 ;
        RECT 84.175 71.015 84.465 71.185 ;
        RECT 84.635 71.015 84.925 71.185 ;
        RECT 85.095 71.015 85.385 71.185 ;
        RECT 85.555 71.015 85.845 71.185 ;
        RECT 86.015 71.015 86.305 71.185 ;
        RECT 86.475 71.015 86.765 71.185 ;
        RECT 86.935 71.015 87.225 71.185 ;
        RECT 87.395 71.015 87.685 71.185 ;
        RECT 87.855 71.015 88.145 71.185 ;
        RECT 88.315 71.015 88.605 71.185 ;
        RECT 88.775 71.015 89.065 71.185 ;
        RECT 89.235 71.015 89.525 71.185 ;
        RECT 89.695 71.015 89.985 71.185 ;
        RECT 90.155 71.015 90.445 71.185 ;
        RECT 90.615 71.015 90.905 71.185 ;
        RECT 91.075 71.015 91.365 71.185 ;
        RECT 91.535 71.015 91.825 71.185 ;
        RECT 91.995 71.015 92.285 71.185 ;
        RECT 92.455 71.015 92.745 71.185 ;
        RECT 92.915 71.015 93.205 71.185 ;
        RECT 93.375 71.015 93.665 71.185 ;
        RECT 93.835 71.015 94.125 71.185 ;
        RECT 94.295 71.015 94.585 71.185 ;
        RECT 94.755 71.015 95.045 71.185 ;
        RECT 95.215 71.015 95.505 71.185 ;
        RECT 95.675 71.015 95.965 71.185 ;
        RECT 96.135 71.015 96.425 71.185 ;
        RECT 96.595 71.015 96.885 71.185 ;
        RECT 97.055 71.015 97.345 71.185 ;
        RECT 97.515 71.015 97.805 71.185 ;
        RECT 97.975 71.015 98.265 71.185 ;
        RECT 98.435 71.015 98.725 71.185 ;
        RECT 98.895 71.015 99.185 71.185 ;
        RECT 99.355 71.015 99.645 71.185 ;
        RECT 99.815 71.015 99.960 71.185 ;
        RECT 16.785 69.925 17.995 71.015 ;
        RECT 18.165 69.925 23.510 71.015 ;
        RECT 23.685 69.925 29.030 71.015 ;
        RECT 29.205 69.925 34.550 71.015 ;
        RECT 34.725 69.925 40.070 71.015 ;
        RECT 40.245 69.925 43.755 71.015 ;
        RECT 16.785 69.215 17.305 69.755 ;
        RECT 17.475 69.385 17.995 69.925 ;
        RECT 18.165 69.235 20.745 69.755 ;
        RECT 20.915 69.405 23.510 69.925 ;
        RECT 23.685 69.235 26.265 69.755 ;
        RECT 26.435 69.405 29.030 69.925 ;
        RECT 29.205 69.235 31.785 69.755 ;
        RECT 31.955 69.405 34.550 69.925 ;
        RECT 34.725 69.235 37.305 69.755 ;
        RECT 37.475 69.405 40.070 69.925 ;
        RECT 40.245 69.235 41.895 69.755 ;
        RECT 42.065 69.405 43.755 69.925 ;
        RECT 44.845 69.850 45.135 71.015 ;
        RECT 45.305 69.925 50.650 71.015 ;
        RECT 50.825 69.925 56.170 71.015 ;
        RECT 56.345 69.925 61.690 71.015 ;
        RECT 61.865 69.925 67.210 71.015 ;
        RECT 67.385 69.925 72.730 71.015 ;
        RECT 45.305 69.235 47.885 69.755 ;
        RECT 48.055 69.405 50.650 69.925 ;
        RECT 50.825 69.235 53.405 69.755 ;
        RECT 53.575 69.405 56.170 69.925 ;
        RECT 56.345 69.235 58.925 69.755 ;
        RECT 59.095 69.405 61.690 69.925 ;
        RECT 61.865 69.235 64.445 69.755 ;
        RECT 64.615 69.405 67.210 69.925 ;
        RECT 67.385 69.235 69.965 69.755 ;
        RECT 70.135 69.405 72.730 69.925 ;
        RECT 72.905 69.850 73.195 71.015 ;
        RECT 73.365 69.925 78.710 71.015 ;
        RECT 78.885 69.925 84.230 71.015 ;
        RECT 84.405 69.925 89.750 71.015 ;
        RECT 89.925 69.925 95.270 71.015 ;
        RECT 95.445 69.925 98.035 71.015 ;
        RECT 73.365 69.235 75.945 69.755 ;
        RECT 76.115 69.405 78.710 69.925 ;
        RECT 78.885 69.235 81.465 69.755 ;
        RECT 81.635 69.405 84.230 69.925 ;
        RECT 84.405 69.235 86.985 69.755 ;
        RECT 87.155 69.405 89.750 69.925 ;
        RECT 89.925 69.235 92.505 69.755 ;
        RECT 92.675 69.405 95.270 69.925 ;
        RECT 95.445 69.235 96.655 69.755 ;
        RECT 96.825 69.405 98.035 69.925 ;
        RECT 98.665 69.925 99.875 71.015 ;
        RECT 98.665 69.385 99.185 69.925 ;
        RECT 16.785 68.465 17.995 69.215 ;
        RECT 18.165 68.465 23.510 69.235 ;
        RECT 23.685 68.465 29.030 69.235 ;
        RECT 29.205 68.465 34.550 69.235 ;
        RECT 34.725 68.465 40.070 69.235 ;
        RECT 40.245 68.465 43.755 69.235 ;
        RECT 44.845 68.465 45.135 69.190 ;
        RECT 45.305 68.465 50.650 69.235 ;
        RECT 50.825 68.465 56.170 69.235 ;
        RECT 56.345 68.465 61.690 69.235 ;
        RECT 61.865 68.465 67.210 69.235 ;
        RECT 67.385 68.465 72.730 69.235 ;
        RECT 72.905 68.465 73.195 69.190 ;
        RECT 73.365 68.465 78.710 69.235 ;
        RECT 78.885 68.465 84.230 69.235 ;
        RECT 84.405 68.465 89.750 69.235 ;
        RECT 89.925 68.465 95.270 69.235 ;
        RECT 95.445 68.465 98.035 69.235 ;
        RECT 99.355 69.215 99.875 69.755 ;
        RECT 98.665 68.465 99.875 69.215 ;
        RECT 16.700 68.295 16.845 68.465 ;
        RECT 17.015 68.295 17.305 68.465 ;
        RECT 17.475 68.295 17.765 68.465 ;
        RECT 17.935 68.295 18.225 68.465 ;
        RECT 18.395 68.295 18.685 68.465 ;
        RECT 18.855 68.295 19.145 68.465 ;
        RECT 19.315 68.295 19.605 68.465 ;
        RECT 19.775 68.295 20.065 68.465 ;
        RECT 20.235 68.295 20.525 68.465 ;
        RECT 20.695 68.295 20.985 68.465 ;
        RECT 21.155 68.295 21.445 68.465 ;
        RECT 21.615 68.295 21.905 68.465 ;
        RECT 22.075 68.295 22.365 68.465 ;
        RECT 22.535 68.295 22.825 68.465 ;
        RECT 22.995 68.295 23.285 68.465 ;
        RECT 23.455 68.295 23.745 68.465 ;
        RECT 23.915 68.295 24.205 68.465 ;
        RECT 24.375 68.295 24.665 68.465 ;
        RECT 24.835 68.295 25.125 68.465 ;
        RECT 25.295 68.295 25.585 68.465 ;
        RECT 25.755 68.295 26.045 68.465 ;
        RECT 26.215 68.295 26.505 68.465 ;
        RECT 26.675 68.295 26.965 68.465 ;
        RECT 27.135 68.295 27.425 68.465 ;
        RECT 27.595 68.295 27.885 68.465 ;
        RECT 28.055 68.295 28.345 68.465 ;
        RECT 28.515 68.295 28.805 68.465 ;
        RECT 28.975 68.295 29.265 68.465 ;
        RECT 29.435 68.295 29.725 68.465 ;
        RECT 29.895 68.295 30.185 68.465 ;
        RECT 30.355 68.295 30.645 68.465 ;
        RECT 30.815 68.295 31.105 68.465 ;
        RECT 31.275 68.295 31.565 68.465 ;
        RECT 31.735 68.295 32.025 68.465 ;
        RECT 32.195 68.295 32.485 68.465 ;
        RECT 32.655 68.295 32.945 68.465 ;
        RECT 33.115 68.295 33.405 68.465 ;
        RECT 33.575 68.295 33.865 68.465 ;
        RECT 34.035 68.295 34.325 68.465 ;
        RECT 34.495 68.295 34.785 68.465 ;
        RECT 34.955 68.295 35.245 68.465 ;
        RECT 35.415 68.295 35.705 68.465 ;
        RECT 35.875 68.295 36.165 68.465 ;
        RECT 36.335 68.295 36.625 68.465 ;
        RECT 36.795 68.295 37.085 68.465 ;
        RECT 37.255 68.295 37.545 68.465 ;
        RECT 37.715 68.295 38.005 68.465 ;
        RECT 38.175 68.295 38.465 68.465 ;
        RECT 38.635 68.295 38.925 68.465 ;
        RECT 39.095 68.295 39.385 68.465 ;
        RECT 39.555 68.295 39.845 68.465 ;
        RECT 40.015 68.295 40.305 68.465 ;
        RECT 40.475 68.295 40.765 68.465 ;
        RECT 40.935 68.295 41.225 68.465 ;
        RECT 41.395 68.295 41.685 68.465 ;
        RECT 41.855 68.295 42.145 68.465 ;
        RECT 42.315 68.295 42.605 68.465 ;
        RECT 42.775 68.295 43.065 68.465 ;
        RECT 43.235 68.295 43.525 68.465 ;
        RECT 43.695 68.295 43.985 68.465 ;
        RECT 44.155 68.295 44.445 68.465 ;
        RECT 44.615 68.295 44.905 68.465 ;
        RECT 45.075 68.295 45.365 68.465 ;
        RECT 45.535 68.295 45.825 68.465 ;
        RECT 45.995 68.295 46.285 68.465 ;
        RECT 46.455 68.295 46.745 68.465 ;
        RECT 46.915 68.295 47.205 68.465 ;
        RECT 47.375 68.295 47.665 68.465 ;
        RECT 47.835 68.295 48.125 68.465 ;
        RECT 48.295 68.295 48.585 68.465 ;
        RECT 48.755 68.295 49.045 68.465 ;
        RECT 49.215 68.295 49.505 68.465 ;
        RECT 49.675 68.295 49.965 68.465 ;
        RECT 50.135 68.295 50.425 68.465 ;
        RECT 50.595 68.295 50.885 68.465 ;
        RECT 51.055 68.295 51.345 68.465 ;
        RECT 51.515 68.295 51.805 68.465 ;
        RECT 51.975 68.295 52.265 68.465 ;
        RECT 52.435 68.295 52.725 68.465 ;
        RECT 52.895 68.295 53.185 68.465 ;
        RECT 53.355 68.295 53.645 68.465 ;
        RECT 53.815 68.295 54.105 68.465 ;
        RECT 54.275 68.295 54.565 68.465 ;
        RECT 54.735 68.295 55.025 68.465 ;
        RECT 55.195 68.295 55.485 68.465 ;
        RECT 55.655 68.295 55.945 68.465 ;
        RECT 56.115 68.295 56.405 68.465 ;
        RECT 56.575 68.295 56.865 68.465 ;
        RECT 57.035 68.295 57.325 68.465 ;
        RECT 57.495 68.295 57.785 68.465 ;
        RECT 57.955 68.295 58.245 68.465 ;
        RECT 58.415 68.295 58.705 68.465 ;
        RECT 58.875 68.295 59.165 68.465 ;
        RECT 59.335 68.295 59.625 68.465 ;
        RECT 59.795 68.295 60.085 68.465 ;
        RECT 60.255 68.295 60.545 68.465 ;
        RECT 60.715 68.295 61.005 68.465 ;
        RECT 61.175 68.295 61.465 68.465 ;
        RECT 61.635 68.295 61.925 68.465 ;
        RECT 62.095 68.295 62.385 68.465 ;
        RECT 62.555 68.295 62.845 68.465 ;
        RECT 63.015 68.295 63.305 68.465 ;
        RECT 63.475 68.295 63.765 68.465 ;
        RECT 63.935 68.295 64.225 68.465 ;
        RECT 64.395 68.295 64.685 68.465 ;
        RECT 64.855 68.295 65.145 68.465 ;
        RECT 65.315 68.295 65.605 68.465 ;
        RECT 65.775 68.295 66.065 68.465 ;
        RECT 66.235 68.295 66.525 68.465 ;
        RECT 66.695 68.295 66.985 68.465 ;
        RECT 67.155 68.295 67.445 68.465 ;
        RECT 67.615 68.295 67.905 68.465 ;
        RECT 68.075 68.295 68.365 68.465 ;
        RECT 68.535 68.295 68.825 68.465 ;
        RECT 68.995 68.295 69.285 68.465 ;
        RECT 69.455 68.295 69.745 68.465 ;
        RECT 69.915 68.295 70.205 68.465 ;
        RECT 70.375 68.295 70.665 68.465 ;
        RECT 70.835 68.295 71.125 68.465 ;
        RECT 71.295 68.295 71.585 68.465 ;
        RECT 71.755 68.295 72.045 68.465 ;
        RECT 72.215 68.295 72.505 68.465 ;
        RECT 72.675 68.295 72.965 68.465 ;
        RECT 73.135 68.295 73.425 68.465 ;
        RECT 73.595 68.295 73.885 68.465 ;
        RECT 74.055 68.295 74.345 68.465 ;
        RECT 74.515 68.295 74.805 68.465 ;
        RECT 74.975 68.295 75.265 68.465 ;
        RECT 75.435 68.295 75.725 68.465 ;
        RECT 75.895 68.295 76.185 68.465 ;
        RECT 76.355 68.295 76.645 68.465 ;
        RECT 76.815 68.295 77.105 68.465 ;
        RECT 77.275 68.295 77.565 68.465 ;
        RECT 77.735 68.295 78.025 68.465 ;
        RECT 78.195 68.295 78.485 68.465 ;
        RECT 78.655 68.295 78.945 68.465 ;
        RECT 79.115 68.295 79.405 68.465 ;
        RECT 79.575 68.295 79.865 68.465 ;
        RECT 80.035 68.295 80.325 68.465 ;
        RECT 80.495 68.295 80.785 68.465 ;
        RECT 80.955 68.295 81.245 68.465 ;
        RECT 81.415 68.295 81.705 68.465 ;
        RECT 81.875 68.295 82.165 68.465 ;
        RECT 82.335 68.295 82.625 68.465 ;
        RECT 82.795 68.295 83.085 68.465 ;
        RECT 83.255 68.295 83.545 68.465 ;
        RECT 83.715 68.295 84.005 68.465 ;
        RECT 84.175 68.295 84.465 68.465 ;
        RECT 84.635 68.295 84.925 68.465 ;
        RECT 85.095 68.295 85.385 68.465 ;
        RECT 85.555 68.295 85.845 68.465 ;
        RECT 86.015 68.295 86.305 68.465 ;
        RECT 86.475 68.295 86.765 68.465 ;
        RECT 86.935 68.295 87.225 68.465 ;
        RECT 87.395 68.295 87.685 68.465 ;
        RECT 87.855 68.295 88.145 68.465 ;
        RECT 88.315 68.295 88.605 68.465 ;
        RECT 88.775 68.295 89.065 68.465 ;
        RECT 89.235 68.295 89.525 68.465 ;
        RECT 89.695 68.295 89.985 68.465 ;
        RECT 90.155 68.295 90.445 68.465 ;
        RECT 90.615 68.295 90.905 68.465 ;
        RECT 91.075 68.295 91.365 68.465 ;
        RECT 91.535 68.295 91.825 68.465 ;
        RECT 91.995 68.295 92.285 68.465 ;
        RECT 92.455 68.295 92.745 68.465 ;
        RECT 92.915 68.295 93.205 68.465 ;
        RECT 93.375 68.295 93.665 68.465 ;
        RECT 93.835 68.295 94.125 68.465 ;
        RECT 94.295 68.295 94.585 68.465 ;
        RECT 94.755 68.295 95.045 68.465 ;
        RECT 95.215 68.295 95.505 68.465 ;
        RECT 95.675 68.295 95.965 68.465 ;
        RECT 96.135 68.295 96.425 68.465 ;
        RECT 96.595 68.295 96.885 68.465 ;
        RECT 97.055 68.295 97.345 68.465 ;
        RECT 97.515 68.295 97.805 68.465 ;
        RECT 97.975 68.295 98.265 68.465 ;
        RECT 98.435 68.295 98.725 68.465 ;
        RECT 98.895 68.295 99.185 68.465 ;
        RECT 99.355 68.295 99.645 68.465 ;
        RECT 99.815 68.295 99.960 68.465 ;
        RECT 16.785 67.545 17.995 68.295 ;
        RECT 16.785 67.005 17.305 67.545 ;
        RECT 18.165 67.525 23.510 68.295 ;
        RECT 23.685 67.525 29.030 68.295 ;
        RECT 29.205 67.525 30.875 68.295 ;
        RECT 31.045 67.570 31.335 68.295 ;
        RECT 31.505 67.525 36.850 68.295 ;
        RECT 37.025 67.525 42.370 68.295 ;
        RECT 42.545 67.525 47.890 68.295 ;
        RECT 48.065 67.525 53.410 68.295 ;
        RECT 53.585 67.525 56.175 68.295 ;
      LAYER li1 ;
        RECT 56.805 67.620 57.065 68.125 ;
      LAYER li1 ;
        RECT 57.245 67.915 57.575 68.295 ;
        RECT 57.755 67.745 57.925 68.125 ;
        RECT 17.475 66.835 17.995 67.375 ;
        RECT 18.165 67.005 20.745 67.525 ;
        RECT 20.915 66.835 23.510 67.355 ;
        RECT 23.685 67.005 26.265 67.525 ;
        RECT 26.435 66.835 29.030 67.355 ;
        RECT 29.205 67.005 29.955 67.525 ;
        RECT 30.125 66.835 30.875 67.355 ;
        RECT 31.505 67.005 34.085 67.525 ;
        RECT 16.785 65.745 17.995 66.835 ;
        RECT 18.165 65.745 23.510 66.835 ;
        RECT 23.685 65.745 29.030 66.835 ;
        RECT 29.205 65.745 30.875 66.835 ;
        RECT 31.045 65.745 31.335 66.910 ;
        RECT 34.255 66.835 36.850 67.355 ;
        RECT 37.025 67.005 39.605 67.525 ;
        RECT 39.775 66.835 42.370 67.355 ;
        RECT 42.545 67.005 45.125 67.525 ;
        RECT 45.295 66.835 47.890 67.355 ;
        RECT 48.065 67.005 50.645 67.525 ;
        RECT 50.815 66.835 53.410 67.355 ;
        RECT 53.585 67.005 54.795 67.525 ;
        RECT 54.965 66.835 56.175 67.355 ;
        RECT 31.505 65.745 36.850 66.835 ;
        RECT 37.025 65.745 42.370 66.835 ;
        RECT 42.545 65.745 47.890 66.835 ;
        RECT 48.065 65.745 53.410 66.835 ;
        RECT 53.585 65.745 56.175 66.835 ;
      LAYER li1 ;
        RECT 56.805 66.820 56.975 67.620 ;
      LAYER li1 ;
        RECT 57.260 67.575 57.925 67.745 ;
        RECT 57.260 67.320 57.430 67.575 ;
        RECT 59.105 67.570 59.395 68.295 ;
        RECT 59.565 67.525 64.910 68.295 ;
        RECT 65.085 67.525 70.430 68.295 ;
        RECT 70.605 67.525 75.950 68.295 ;
        RECT 76.125 67.525 81.470 68.295 ;
        RECT 81.645 67.525 86.990 68.295 ;
        RECT 87.165 67.570 87.455 68.295 ;
        RECT 87.625 67.525 92.970 68.295 ;
        RECT 93.145 67.525 98.490 68.295 ;
        RECT 98.665 67.545 99.875 68.295 ;
        RECT 57.145 66.990 57.430 67.320 ;
      LAYER li1 ;
        RECT 57.665 67.025 57.995 67.395 ;
      LAYER li1 ;
        RECT 59.565 67.005 62.145 67.525 ;
        RECT 57.260 66.845 57.430 66.990 ;
      LAYER li1 ;
        RECT 56.805 65.915 57.075 66.820 ;
      LAYER li1 ;
        RECT 57.260 66.675 57.925 66.845 ;
        RECT 57.245 65.745 57.575 66.505 ;
        RECT 57.755 65.915 57.925 66.675 ;
        RECT 59.105 65.745 59.395 66.910 ;
        RECT 62.315 66.835 64.910 67.355 ;
        RECT 65.085 67.005 67.665 67.525 ;
        RECT 67.835 66.835 70.430 67.355 ;
        RECT 70.605 67.005 73.185 67.525 ;
        RECT 73.355 66.835 75.950 67.355 ;
        RECT 76.125 67.005 78.705 67.525 ;
        RECT 78.875 66.835 81.470 67.355 ;
        RECT 81.645 67.005 84.225 67.525 ;
        RECT 84.395 66.835 86.990 67.355 ;
        RECT 87.625 67.005 90.205 67.525 ;
        RECT 59.565 65.745 64.910 66.835 ;
        RECT 65.085 65.745 70.430 66.835 ;
        RECT 70.605 65.745 75.950 66.835 ;
        RECT 76.125 65.745 81.470 66.835 ;
        RECT 81.645 65.745 86.990 66.835 ;
        RECT 87.165 65.745 87.455 66.910 ;
        RECT 90.375 66.835 92.970 67.355 ;
        RECT 93.145 67.005 95.725 67.525 ;
        RECT 95.895 66.835 98.490 67.355 ;
        RECT 87.625 65.745 92.970 66.835 ;
        RECT 93.145 65.745 98.490 66.835 ;
        RECT 98.665 66.835 99.185 67.375 ;
        RECT 99.355 67.005 99.875 67.545 ;
        RECT 98.665 65.745 99.875 66.835 ;
        RECT 16.700 65.575 16.845 65.745 ;
        RECT 17.015 65.575 17.305 65.745 ;
        RECT 17.475 65.575 17.765 65.745 ;
        RECT 17.935 65.575 18.225 65.745 ;
        RECT 18.395 65.575 18.685 65.745 ;
        RECT 18.855 65.575 19.145 65.745 ;
        RECT 19.315 65.575 19.605 65.745 ;
        RECT 19.775 65.575 20.065 65.745 ;
        RECT 20.235 65.575 20.525 65.745 ;
        RECT 20.695 65.575 20.985 65.745 ;
        RECT 21.155 65.575 21.445 65.745 ;
        RECT 21.615 65.575 21.905 65.745 ;
        RECT 22.075 65.575 22.365 65.745 ;
        RECT 22.535 65.575 22.825 65.745 ;
        RECT 22.995 65.575 23.285 65.745 ;
        RECT 23.455 65.575 23.745 65.745 ;
        RECT 23.915 65.575 24.205 65.745 ;
        RECT 24.375 65.575 24.665 65.745 ;
        RECT 24.835 65.575 25.125 65.745 ;
        RECT 25.295 65.575 25.585 65.745 ;
        RECT 25.755 65.575 26.045 65.745 ;
        RECT 26.215 65.575 26.505 65.745 ;
        RECT 26.675 65.575 26.965 65.745 ;
        RECT 27.135 65.575 27.425 65.745 ;
        RECT 27.595 65.575 27.885 65.745 ;
        RECT 28.055 65.575 28.345 65.745 ;
        RECT 28.515 65.575 28.805 65.745 ;
        RECT 28.975 65.575 29.265 65.745 ;
        RECT 29.435 65.575 29.725 65.745 ;
        RECT 29.895 65.575 30.185 65.745 ;
        RECT 30.355 65.575 30.645 65.745 ;
        RECT 30.815 65.575 31.105 65.745 ;
        RECT 31.275 65.575 31.565 65.745 ;
        RECT 31.735 65.575 32.025 65.745 ;
        RECT 32.195 65.575 32.485 65.745 ;
        RECT 32.655 65.575 32.945 65.745 ;
        RECT 33.115 65.575 33.405 65.745 ;
        RECT 33.575 65.575 33.865 65.745 ;
        RECT 34.035 65.575 34.325 65.745 ;
        RECT 34.495 65.575 34.785 65.745 ;
        RECT 34.955 65.575 35.245 65.745 ;
        RECT 35.415 65.575 35.705 65.745 ;
        RECT 35.875 65.575 36.165 65.745 ;
        RECT 36.335 65.575 36.625 65.745 ;
        RECT 36.795 65.575 37.085 65.745 ;
        RECT 37.255 65.575 37.545 65.745 ;
        RECT 37.715 65.575 38.005 65.745 ;
        RECT 38.175 65.575 38.465 65.745 ;
        RECT 38.635 65.575 38.925 65.745 ;
        RECT 39.095 65.575 39.385 65.745 ;
        RECT 39.555 65.575 39.845 65.745 ;
        RECT 40.015 65.575 40.305 65.745 ;
        RECT 40.475 65.575 40.765 65.745 ;
        RECT 40.935 65.575 41.225 65.745 ;
        RECT 41.395 65.575 41.685 65.745 ;
        RECT 41.855 65.575 42.145 65.745 ;
        RECT 42.315 65.575 42.605 65.745 ;
        RECT 42.775 65.575 43.065 65.745 ;
        RECT 43.235 65.575 43.525 65.745 ;
        RECT 43.695 65.575 43.985 65.745 ;
        RECT 44.155 65.575 44.445 65.745 ;
        RECT 44.615 65.575 44.905 65.745 ;
        RECT 45.075 65.575 45.365 65.745 ;
        RECT 45.535 65.575 45.825 65.745 ;
        RECT 45.995 65.575 46.285 65.745 ;
        RECT 46.455 65.575 46.745 65.745 ;
        RECT 46.915 65.575 47.205 65.745 ;
        RECT 47.375 65.575 47.665 65.745 ;
        RECT 47.835 65.575 48.125 65.745 ;
        RECT 48.295 65.575 48.585 65.745 ;
        RECT 48.755 65.575 49.045 65.745 ;
        RECT 49.215 65.575 49.505 65.745 ;
        RECT 49.675 65.575 49.965 65.745 ;
        RECT 50.135 65.575 50.425 65.745 ;
        RECT 50.595 65.575 50.885 65.745 ;
        RECT 51.055 65.575 51.345 65.745 ;
        RECT 51.515 65.575 51.805 65.745 ;
        RECT 51.975 65.575 52.265 65.745 ;
        RECT 52.435 65.575 52.725 65.745 ;
        RECT 52.895 65.575 53.185 65.745 ;
        RECT 53.355 65.575 53.645 65.745 ;
        RECT 53.815 65.575 54.105 65.745 ;
        RECT 54.275 65.575 54.565 65.745 ;
        RECT 54.735 65.575 55.025 65.745 ;
        RECT 55.195 65.575 55.485 65.745 ;
        RECT 55.655 65.575 55.945 65.745 ;
        RECT 56.115 65.575 56.405 65.745 ;
        RECT 56.575 65.575 56.865 65.745 ;
        RECT 57.035 65.575 57.325 65.745 ;
        RECT 57.495 65.575 57.785 65.745 ;
        RECT 57.955 65.575 58.245 65.745 ;
        RECT 58.415 65.575 58.705 65.745 ;
        RECT 58.875 65.575 59.165 65.745 ;
        RECT 59.335 65.575 59.625 65.745 ;
        RECT 59.795 65.575 60.085 65.745 ;
        RECT 60.255 65.575 60.545 65.745 ;
        RECT 60.715 65.575 61.005 65.745 ;
        RECT 61.175 65.575 61.465 65.745 ;
        RECT 61.635 65.575 61.925 65.745 ;
        RECT 62.095 65.575 62.385 65.745 ;
        RECT 62.555 65.575 62.845 65.745 ;
        RECT 63.015 65.575 63.305 65.745 ;
        RECT 63.475 65.575 63.765 65.745 ;
        RECT 63.935 65.575 64.225 65.745 ;
        RECT 64.395 65.575 64.685 65.745 ;
        RECT 64.855 65.575 65.145 65.745 ;
        RECT 65.315 65.575 65.605 65.745 ;
        RECT 65.775 65.575 66.065 65.745 ;
        RECT 66.235 65.575 66.525 65.745 ;
        RECT 66.695 65.575 66.985 65.745 ;
        RECT 67.155 65.575 67.445 65.745 ;
        RECT 67.615 65.575 67.905 65.745 ;
        RECT 68.075 65.575 68.365 65.745 ;
        RECT 68.535 65.575 68.825 65.745 ;
        RECT 68.995 65.575 69.285 65.745 ;
        RECT 69.455 65.575 69.745 65.745 ;
        RECT 69.915 65.575 70.205 65.745 ;
        RECT 70.375 65.575 70.665 65.745 ;
        RECT 70.835 65.575 71.125 65.745 ;
        RECT 71.295 65.575 71.585 65.745 ;
        RECT 71.755 65.575 72.045 65.745 ;
        RECT 72.215 65.575 72.505 65.745 ;
        RECT 72.675 65.575 72.965 65.745 ;
        RECT 73.135 65.575 73.425 65.745 ;
        RECT 73.595 65.575 73.885 65.745 ;
        RECT 74.055 65.575 74.345 65.745 ;
        RECT 74.515 65.575 74.805 65.745 ;
        RECT 74.975 65.575 75.265 65.745 ;
        RECT 75.435 65.575 75.725 65.745 ;
        RECT 75.895 65.575 76.185 65.745 ;
        RECT 76.355 65.575 76.645 65.745 ;
        RECT 76.815 65.575 77.105 65.745 ;
        RECT 77.275 65.575 77.565 65.745 ;
        RECT 77.735 65.575 78.025 65.745 ;
        RECT 78.195 65.575 78.485 65.745 ;
        RECT 78.655 65.575 78.945 65.745 ;
        RECT 79.115 65.575 79.405 65.745 ;
        RECT 79.575 65.575 79.865 65.745 ;
        RECT 80.035 65.575 80.325 65.745 ;
        RECT 80.495 65.575 80.785 65.745 ;
        RECT 80.955 65.575 81.245 65.745 ;
        RECT 81.415 65.575 81.705 65.745 ;
        RECT 81.875 65.575 82.165 65.745 ;
        RECT 82.335 65.575 82.625 65.745 ;
        RECT 82.795 65.575 83.085 65.745 ;
        RECT 83.255 65.575 83.545 65.745 ;
        RECT 83.715 65.575 84.005 65.745 ;
        RECT 84.175 65.575 84.465 65.745 ;
        RECT 84.635 65.575 84.925 65.745 ;
        RECT 85.095 65.575 85.385 65.745 ;
        RECT 85.555 65.575 85.845 65.745 ;
        RECT 86.015 65.575 86.305 65.745 ;
        RECT 86.475 65.575 86.765 65.745 ;
        RECT 86.935 65.575 87.225 65.745 ;
        RECT 87.395 65.575 87.685 65.745 ;
        RECT 87.855 65.575 88.145 65.745 ;
        RECT 88.315 65.575 88.605 65.745 ;
        RECT 88.775 65.575 89.065 65.745 ;
        RECT 89.235 65.575 89.525 65.745 ;
        RECT 89.695 65.575 89.985 65.745 ;
        RECT 90.155 65.575 90.445 65.745 ;
        RECT 90.615 65.575 90.905 65.745 ;
        RECT 91.075 65.575 91.365 65.745 ;
        RECT 91.535 65.575 91.825 65.745 ;
        RECT 91.995 65.575 92.285 65.745 ;
        RECT 92.455 65.575 92.745 65.745 ;
        RECT 92.915 65.575 93.205 65.745 ;
        RECT 93.375 65.575 93.665 65.745 ;
        RECT 93.835 65.575 94.125 65.745 ;
        RECT 94.295 65.575 94.585 65.745 ;
        RECT 94.755 65.575 95.045 65.745 ;
        RECT 95.215 65.575 95.505 65.745 ;
        RECT 95.675 65.575 95.965 65.745 ;
        RECT 96.135 65.575 96.425 65.745 ;
        RECT 96.595 65.575 96.885 65.745 ;
        RECT 97.055 65.575 97.345 65.745 ;
        RECT 97.515 65.575 97.805 65.745 ;
        RECT 97.975 65.575 98.265 65.745 ;
        RECT 98.435 65.575 98.725 65.745 ;
        RECT 98.895 65.575 99.185 65.745 ;
        RECT 99.355 65.575 99.645 65.745 ;
        RECT 99.815 65.575 99.960 65.745 ;
        RECT 16.785 64.485 17.995 65.575 ;
        RECT 18.165 64.485 23.510 65.575 ;
        RECT 23.685 64.485 29.030 65.575 ;
        RECT 29.205 64.485 34.550 65.575 ;
        RECT 34.725 64.485 40.070 65.575 ;
        RECT 40.245 64.485 43.755 65.575 ;
        RECT 16.785 63.775 17.305 64.315 ;
        RECT 17.475 63.945 17.995 64.485 ;
        RECT 18.165 63.795 20.745 64.315 ;
        RECT 20.915 63.965 23.510 64.485 ;
        RECT 23.685 63.795 26.265 64.315 ;
        RECT 26.435 63.965 29.030 64.485 ;
        RECT 29.205 63.795 31.785 64.315 ;
        RECT 31.955 63.965 34.550 64.485 ;
        RECT 34.725 63.795 37.305 64.315 ;
        RECT 37.475 63.965 40.070 64.485 ;
        RECT 40.245 63.795 41.895 64.315 ;
        RECT 42.065 63.965 43.755 64.485 ;
        RECT 44.845 64.410 45.135 65.575 ;
        RECT 45.305 64.485 50.650 65.575 ;
        RECT 50.825 64.485 56.170 65.575 ;
        RECT 56.345 64.485 59.855 65.575 ;
        RECT 60.575 64.905 60.745 65.405 ;
        RECT 60.915 65.075 61.245 65.575 ;
        RECT 60.575 64.735 61.240 64.905 ;
        RECT 45.305 63.795 47.885 64.315 ;
        RECT 48.055 63.965 50.650 64.485 ;
        RECT 50.825 63.795 53.405 64.315 ;
        RECT 53.575 63.965 56.170 64.485 ;
        RECT 56.345 63.795 57.995 64.315 ;
        RECT 58.165 63.965 59.855 64.485 ;
      LAYER li1 ;
        RECT 60.490 63.915 60.840 64.565 ;
      LAYER li1 ;
        RECT 16.785 63.025 17.995 63.775 ;
        RECT 18.165 63.025 23.510 63.795 ;
        RECT 23.685 63.025 29.030 63.795 ;
        RECT 29.205 63.025 34.550 63.795 ;
        RECT 34.725 63.025 40.070 63.795 ;
        RECT 40.245 63.025 43.755 63.795 ;
        RECT 44.845 63.025 45.135 63.750 ;
        RECT 45.305 63.025 50.650 63.795 ;
        RECT 50.825 63.025 56.170 63.795 ;
        RECT 56.345 63.025 59.855 63.795 ;
        RECT 61.010 63.745 61.240 64.735 ;
        RECT 60.575 63.575 61.240 63.745 ;
        RECT 60.575 63.285 60.745 63.575 ;
        RECT 60.915 63.025 61.245 63.405 ;
        RECT 61.415 63.285 61.640 65.405 ;
        RECT 61.840 65.115 62.105 65.575 ;
        RECT 62.290 65.005 62.525 65.380 ;
        RECT 62.770 65.130 63.840 65.300 ;
      LAYER li1 ;
        RECT 61.840 64.005 62.120 64.605 ;
      LAYER li1 ;
        RECT 61.855 63.025 62.105 63.485 ;
        RECT 62.290 63.475 62.460 65.005 ;
        RECT 62.630 63.975 62.870 64.845 ;
        RECT 63.060 64.595 63.500 64.950 ;
        RECT 63.670 64.515 63.840 65.130 ;
        RECT 64.010 64.775 64.180 65.575 ;
        RECT 64.350 65.075 64.600 65.405 ;
        RECT 64.825 65.105 65.710 65.275 ;
        RECT 63.670 64.425 64.180 64.515 ;
        RECT 63.380 64.255 64.180 64.425 ;
        RECT 62.630 63.645 63.210 63.975 ;
        RECT 63.380 63.475 63.550 64.255 ;
        RECT 64.010 64.185 64.180 64.255 ;
        RECT 63.720 64.005 63.890 64.035 ;
        RECT 64.350 64.005 64.520 65.075 ;
        RECT 64.690 64.185 64.880 64.905 ;
        RECT 65.050 64.515 65.370 64.845 ;
        RECT 63.720 63.705 64.520 64.005 ;
        RECT 65.050 63.975 65.240 64.515 ;
        RECT 62.290 63.305 62.620 63.475 ;
        RECT 62.800 63.305 63.550 63.475 ;
        RECT 63.800 63.025 64.170 63.525 ;
        RECT 64.350 63.475 64.520 63.705 ;
        RECT 64.690 63.645 65.240 63.975 ;
        RECT 65.540 64.185 65.710 65.105 ;
        RECT 65.890 65.075 66.105 65.575 ;
        RECT 66.570 64.770 66.740 65.395 ;
        RECT 67.025 64.795 67.205 65.575 ;
        RECT 65.880 64.610 66.740 64.770 ;
        RECT 67.900 64.745 68.070 65.575 ;
        RECT 68.740 64.745 68.910 65.575 ;
        RECT 65.880 64.440 66.990 64.610 ;
        RECT 69.225 64.485 72.735 65.575 ;
        RECT 66.820 64.185 66.990 64.440 ;
        RECT 65.540 64.015 66.630 64.185 ;
        RECT 66.820 64.015 68.640 64.185 ;
        RECT 65.540 63.475 65.710 64.015 ;
        RECT 66.820 63.845 66.990 64.015 ;
        RECT 66.490 63.675 66.990 63.845 ;
        RECT 69.225 63.795 70.875 64.315 ;
        RECT 71.045 63.965 72.735 64.485 ;
        RECT 72.905 64.410 73.195 65.575 ;
        RECT 73.365 64.485 78.710 65.575 ;
        RECT 78.885 64.485 84.230 65.575 ;
        RECT 84.405 64.485 89.750 65.575 ;
        RECT 89.925 64.485 95.270 65.575 ;
        RECT 95.445 64.485 98.035 65.575 ;
        RECT 73.365 63.795 75.945 64.315 ;
        RECT 76.115 63.965 78.710 64.485 ;
        RECT 78.885 63.795 81.465 64.315 ;
        RECT 81.635 63.965 84.230 64.485 ;
        RECT 84.405 63.795 86.985 64.315 ;
        RECT 87.155 63.965 89.750 64.485 ;
        RECT 89.925 63.795 92.505 64.315 ;
        RECT 92.675 63.965 95.270 64.485 ;
        RECT 95.445 63.795 96.655 64.315 ;
        RECT 96.825 63.965 98.035 64.485 ;
        RECT 98.665 64.485 99.875 65.575 ;
        RECT 98.665 63.945 99.185 64.485 ;
        RECT 64.350 63.305 64.810 63.475 ;
        RECT 65.040 63.305 65.710 63.475 ;
        RECT 66.025 63.025 66.195 63.555 ;
        RECT 66.490 63.235 66.850 63.675 ;
        RECT 67.025 63.025 67.195 63.505 ;
        RECT 67.895 63.025 68.065 63.500 ;
        RECT 68.745 63.025 68.915 63.500 ;
        RECT 69.225 63.025 72.735 63.795 ;
        RECT 72.905 63.025 73.195 63.750 ;
        RECT 73.365 63.025 78.710 63.795 ;
        RECT 78.885 63.025 84.230 63.795 ;
        RECT 84.405 63.025 89.750 63.795 ;
        RECT 89.925 63.025 95.270 63.795 ;
        RECT 95.445 63.025 98.035 63.795 ;
        RECT 99.355 63.775 99.875 64.315 ;
        RECT 98.665 63.025 99.875 63.775 ;
        RECT 16.700 62.855 16.845 63.025 ;
        RECT 17.015 62.855 17.305 63.025 ;
        RECT 17.475 62.855 17.765 63.025 ;
        RECT 17.935 62.855 18.225 63.025 ;
        RECT 18.395 62.855 18.685 63.025 ;
        RECT 18.855 62.855 19.145 63.025 ;
        RECT 19.315 62.855 19.605 63.025 ;
        RECT 19.775 62.855 20.065 63.025 ;
        RECT 20.235 62.855 20.525 63.025 ;
        RECT 20.695 62.855 20.985 63.025 ;
        RECT 21.155 62.855 21.445 63.025 ;
        RECT 21.615 62.855 21.905 63.025 ;
        RECT 22.075 62.855 22.365 63.025 ;
        RECT 22.535 62.855 22.825 63.025 ;
        RECT 22.995 62.855 23.285 63.025 ;
        RECT 23.455 62.855 23.745 63.025 ;
        RECT 23.915 62.855 24.205 63.025 ;
        RECT 24.375 62.855 24.665 63.025 ;
        RECT 24.835 62.855 25.125 63.025 ;
        RECT 25.295 62.855 25.585 63.025 ;
        RECT 25.755 62.855 26.045 63.025 ;
        RECT 26.215 62.855 26.505 63.025 ;
        RECT 26.675 62.855 26.965 63.025 ;
        RECT 27.135 62.855 27.425 63.025 ;
        RECT 27.595 62.855 27.885 63.025 ;
        RECT 28.055 62.855 28.345 63.025 ;
        RECT 28.515 62.855 28.805 63.025 ;
        RECT 28.975 62.855 29.265 63.025 ;
        RECT 29.435 62.855 29.725 63.025 ;
        RECT 29.895 62.855 30.185 63.025 ;
        RECT 30.355 62.855 30.645 63.025 ;
        RECT 30.815 62.855 31.105 63.025 ;
        RECT 31.275 62.855 31.565 63.025 ;
        RECT 31.735 62.855 32.025 63.025 ;
        RECT 32.195 62.855 32.485 63.025 ;
        RECT 32.655 62.855 32.945 63.025 ;
        RECT 33.115 62.855 33.405 63.025 ;
        RECT 33.575 62.855 33.865 63.025 ;
        RECT 34.035 62.855 34.325 63.025 ;
        RECT 34.495 62.855 34.785 63.025 ;
        RECT 34.955 62.855 35.245 63.025 ;
        RECT 35.415 62.855 35.705 63.025 ;
        RECT 35.875 62.855 36.165 63.025 ;
        RECT 36.335 62.855 36.625 63.025 ;
        RECT 36.795 62.855 37.085 63.025 ;
        RECT 37.255 62.855 37.545 63.025 ;
        RECT 37.715 62.855 38.005 63.025 ;
        RECT 38.175 62.855 38.465 63.025 ;
        RECT 38.635 62.855 38.925 63.025 ;
        RECT 39.095 62.855 39.385 63.025 ;
        RECT 39.555 62.855 39.845 63.025 ;
        RECT 40.015 62.855 40.305 63.025 ;
        RECT 40.475 62.855 40.765 63.025 ;
        RECT 40.935 62.855 41.225 63.025 ;
        RECT 41.395 62.855 41.685 63.025 ;
        RECT 41.855 62.855 42.145 63.025 ;
        RECT 42.315 62.855 42.605 63.025 ;
        RECT 42.775 62.855 43.065 63.025 ;
        RECT 43.235 62.855 43.525 63.025 ;
        RECT 43.695 62.855 43.985 63.025 ;
        RECT 44.155 62.855 44.445 63.025 ;
        RECT 44.615 62.855 44.905 63.025 ;
        RECT 45.075 62.855 45.365 63.025 ;
        RECT 45.535 62.855 45.825 63.025 ;
        RECT 45.995 62.855 46.285 63.025 ;
        RECT 46.455 62.855 46.745 63.025 ;
        RECT 46.915 62.855 47.205 63.025 ;
        RECT 47.375 62.855 47.665 63.025 ;
        RECT 47.835 62.855 48.125 63.025 ;
        RECT 48.295 62.855 48.585 63.025 ;
        RECT 48.755 62.855 49.045 63.025 ;
        RECT 49.215 62.855 49.505 63.025 ;
        RECT 49.675 62.855 49.965 63.025 ;
        RECT 50.135 62.855 50.425 63.025 ;
        RECT 50.595 62.855 50.885 63.025 ;
        RECT 51.055 62.855 51.345 63.025 ;
        RECT 51.515 62.855 51.805 63.025 ;
        RECT 51.975 62.855 52.265 63.025 ;
        RECT 52.435 62.855 52.725 63.025 ;
        RECT 52.895 62.855 53.185 63.025 ;
        RECT 53.355 62.855 53.645 63.025 ;
        RECT 53.815 62.855 54.105 63.025 ;
        RECT 54.275 62.855 54.565 63.025 ;
        RECT 54.735 62.855 55.025 63.025 ;
        RECT 55.195 62.855 55.485 63.025 ;
        RECT 55.655 62.855 55.945 63.025 ;
        RECT 56.115 62.855 56.405 63.025 ;
        RECT 56.575 62.855 56.865 63.025 ;
        RECT 57.035 62.855 57.325 63.025 ;
        RECT 57.495 62.855 57.785 63.025 ;
        RECT 57.955 62.855 58.245 63.025 ;
        RECT 58.415 62.855 58.705 63.025 ;
        RECT 58.875 62.855 59.165 63.025 ;
        RECT 59.335 62.855 59.625 63.025 ;
        RECT 59.795 62.855 60.085 63.025 ;
        RECT 60.255 62.855 60.545 63.025 ;
        RECT 60.715 62.855 61.005 63.025 ;
        RECT 61.175 62.855 61.465 63.025 ;
        RECT 61.635 62.855 61.925 63.025 ;
        RECT 62.095 62.855 62.385 63.025 ;
        RECT 62.555 62.855 62.845 63.025 ;
        RECT 63.015 62.855 63.305 63.025 ;
        RECT 63.475 62.855 63.765 63.025 ;
        RECT 63.935 62.855 64.225 63.025 ;
        RECT 64.395 62.855 64.685 63.025 ;
        RECT 64.855 62.855 65.145 63.025 ;
        RECT 65.315 62.855 65.605 63.025 ;
        RECT 65.775 62.855 66.065 63.025 ;
        RECT 66.235 62.855 66.525 63.025 ;
        RECT 66.695 62.855 66.985 63.025 ;
        RECT 67.155 62.855 67.445 63.025 ;
        RECT 67.615 62.855 67.905 63.025 ;
        RECT 68.075 62.855 68.365 63.025 ;
        RECT 68.535 62.855 68.825 63.025 ;
        RECT 68.995 62.855 69.285 63.025 ;
        RECT 69.455 62.855 69.745 63.025 ;
        RECT 69.915 62.855 70.205 63.025 ;
        RECT 70.375 62.855 70.665 63.025 ;
        RECT 70.835 62.855 71.125 63.025 ;
        RECT 71.295 62.855 71.585 63.025 ;
        RECT 71.755 62.855 72.045 63.025 ;
        RECT 72.215 62.855 72.505 63.025 ;
        RECT 72.675 62.855 72.965 63.025 ;
        RECT 73.135 62.855 73.425 63.025 ;
        RECT 73.595 62.855 73.885 63.025 ;
        RECT 74.055 62.855 74.345 63.025 ;
        RECT 74.515 62.855 74.805 63.025 ;
        RECT 74.975 62.855 75.265 63.025 ;
        RECT 75.435 62.855 75.725 63.025 ;
        RECT 75.895 62.855 76.185 63.025 ;
        RECT 76.355 62.855 76.645 63.025 ;
        RECT 76.815 62.855 77.105 63.025 ;
        RECT 77.275 62.855 77.565 63.025 ;
        RECT 77.735 62.855 78.025 63.025 ;
        RECT 78.195 62.855 78.485 63.025 ;
        RECT 78.655 62.855 78.945 63.025 ;
        RECT 79.115 62.855 79.405 63.025 ;
        RECT 79.575 62.855 79.865 63.025 ;
        RECT 80.035 62.855 80.325 63.025 ;
        RECT 80.495 62.855 80.785 63.025 ;
        RECT 80.955 62.855 81.245 63.025 ;
        RECT 81.415 62.855 81.705 63.025 ;
        RECT 81.875 62.855 82.165 63.025 ;
        RECT 82.335 62.855 82.625 63.025 ;
        RECT 82.795 62.855 83.085 63.025 ;
        RECT 83.255 62.855 83.545 63.025 ;
        RECT 83.715 62.855 84.005 63.025 ;
        RECT 84.175 62.855 84.465 63.025 ;
        RECT 84.635 62.855 84.925 63.025 ;
        RECT 85.095 62.855 85.385 63.025 ;
        RECT 85.555 62.855 85.845 63.025 ;
        RECT 86.015 62.855 86.305 63.025 ;
        RECT 86.475 62.855 86.765 63.025 ;
        RECT 86.935 62.855 87.225 63.025 ;
        RECT 87.395 62.855 87.685 63.025 ;
        RECT 87.855 62.855 88.145 63.025 ;
        RECT 88.315 62.855 88.605 63.025 ;
        RECT 88.775 62.855 89.065 63.025 ;
        RECT 89.235 62.855 89.525 63.025 ;
        RECT 89.695 62.855 89.985 63.025 ;
        RECT 90.155 62.855 90.445 63.025 ;
        RECT 90.615 62.855 90.905 63.025 ;
        RECT 91.075 62.855 91.365 63.025 ;
        RECT 91.535 62.855 91.825 63.025 ;
        RECT 91.995 62.855 92.285 63.025 ;
        RECT 92.455 62.855 92.745 63.025 ;
        RECT 92.915 62.855 93.205 63.025 ;
        RECT 93.375 62.855 93.665 63.025 ;
        RECT 93.835 62.855 94.125 63.025 ;
        RECT 94.295 62.855 94.585 63.025 ;
        RECT 94.755 62.855 95.045 63.025 ;
        RECT 95.215 62.855 95.505 63.025 ;
        RECT 95.675 62.855 95.965 63.025 ;
        RECT 96.135 62.855 96.425 63.025 ;
        RECT 96.595 62.855 96.885 63.025 ;
        RECT 97.055 62.855 97.345 63.025 ;
        RECT 97.515 62.855 97.805 63.025 ;
        RECT 97.975 62.855 98.265 63.025 ;
        RECT 98.435 62.855 98.725 63.025 ;
        RECT 98.895 62.855 99.185 63.025 ;
        RECT 99.355 62.855 99.645 63.025 ;
        RECT 99.815 62.855 99.960 63.025 ;
        RECT 16.785 62.105 17.995 62.855 ;
        RECT 18.165 62.105 19.375 62.855 ;
        RECT 16.785 61.565 17.305 62.105 ;
        RECT 17.475 61.395 17.995 61.935 ;
        RECT 18.165 61.565 18.685 62.105 ;
        RECT 18.855 61.395 19.375 61.935 ;
        RECT 16.785 60.305 17.995 61.395 ;
        RECT 18.165 60.305 19.375 61.395 ;
      LAYER li1 ;
        RECT 19.545 61.200 20.065 62.685 ;
      LAYER li1 ;
        RECT 20.235 62.195 20.575 62.855 ;
        RECT 20.925 62.085 26.270 62.855 ;
        RECT 26.445 62.085 29.955 62.855 ;
        RECT 31.045 62.130 31.335 62.855 ;
        RECT 31.505 62.085 36.850 62.855 ;
        RECT 37.025 62.085 40.535 62.855 ;
        RECT 40.795 62.305 40.965 62.595 ;
        RECT 41.135 62.475 41.465 62.855 ;
        RECT 40.795 62.135 41.460 62.305 ;
        RECT 20.925 61.565 23.505 62.085 ;
        RECT 23.675 61.395 26.270 61.915 ;
        RECT 26.445 61.565 28.095 62.085 ;
        RECT 28.265 61.395 29.955 61.915 ;
        RECT 31.505 61.565 34.085 62.085 ;
        RECT 19.735 60.305 20.065 61.030 ;
        RECT 20.925 60.305 26.270 61.395 ;
        RECT 26.445 60.305 29.955 61.395 ;
        RECT 31.045 60.305 31.335 61.470 ;
        RECT 34.255 61.395 36.850 61.915 ;
        RECT 37.025 61.565 38.675 62.085 ;
        RECT 38.845 61.395 40.535 61.915 ;
        RECT 31.505 60.305 36.850 61.395 ;
        RECT 37.025 60.305 40.535 61.395 ;
      LAYER li1 ;
        RECT 40.710 61.315 41.060 61.965 ;
      LAYER li1 ;
        RECT 41.230 61.145 41.460 62.135 ;
        RECT 40.795 60.975 41.460 61.145 ;
        RECT 40.795 60.475 40.965 60.975 ;
        RECT 41.135 60.305 41.465 60.805 ;
        RECT 41.635 60.475 41.860 62.595 ;
        RECT 42.075 62.395 42.325 62.855 ;
        RECT 42.510 62.405 42.840 62.575 ;
        RECT 43.020 62.405 43.770 62.575 ;
      LAYER li1 ;
        RECT 42.060 61.275 42.340 61.875 ;
      LAYER li1 ;
        RECT 42.510 60.875 42.680 62.405 ;
        RECT 42.850 61.905 43.430 62.235 ;
        RECT 42.850 61.035 43.090 61.905 ;
        RECT 43.600 61.625 43.770 62.405 ;
        RECT 44.020 62.355 44.390 62.855 ;
        RECT 44.570 62.405 45.030 62.575 ;
        RECT 45.260 62.405 45.930 62.575 ;
        RECT 44.570 62.175 44.740 62.405 ;
        RECT 43.940 61.875 44.740 62.175 ;
        RECT 44.910 61.905 45.460 62.235 ;
        RECT 43.940 61.845 44.110 61.875 ;
        RECT 44.230 61.625 44.400 61.695 ;
        RECT 43.600 61.455 44.400 61.625 ;
        RECT 43.890 61.365 44.400 61.455 ;
        RECT 43.280 60.930 43.720 61.285 ;
        RECT 42.060 60.305 42.325 60.765 ;
        RECT 42.510 60.500 42.745 60.875 ;
        RECT 43.890 60.750 44.060 61.365 ;
        RECT 42.990 60.580 44.060 60.750 ;
        RECT 44.230 60.305 44.400 61.105 ;
        RECT 44.570 60.805 44.740 61.875 ;
        RECT 44.910 60.975 45.100 61.695 ;
        RECT 45.270 61.365 45.460 61.905 ;
        RECT 45.760 61.865 45.930 62.405 ;
        RECT 46.245 62.325 46.415 62.855 ;
        RECT 46.710 62.205 47.070 62.645 ;
        RECT 47.245 62.375 47.415 62.855 ;
        RECT 48.115 62.380 48.285 62.855 ;
        RECT 48.965 62.380 49.135 62.855 ;
        RECT 46.710 62.035 47.210 62.205 ;
        RECT 47.040 61.865 47.210 62.035 ;
        RECT 49.445 62.085 54.790 62.855 ;
        RECT 54.965 62.085 58.475 62.855 ;
        RECT 59.105 62.130 59.395 62.855 ;
        RECT 60.115 62.305 60.285 62.685 ;
        RECT 60.500 62.475 60.830 62.855 ;
        RECT 60.115 62.135 60.830 62.305 ;
        RECT 45.760 61.695 46.850 61.865 ;
        RECT 47.040 61.695 48.860 61.865 ;
        RECT 45.270 61.035 45.590 61.365 ;
        RECT 44.570 60.475 44.820 60.805 ;
        RECT 45.760 60.775 45.930 61.695 ;
        RECT 47.040 61.440 47.210 61.695 ;
        RECT 49.445 61.565 52.025 62.085 ;
        RECT 46.100 61.270 47.210 61.440 ;
        RECT 52.195 61.395 54.790 61.915 ;
        RECT 54.965 61.565 56.615 62.085 ;
        RECT 56.785 61.395 58.475 61.915 ;
      LAYER li1 ;
        RECT 60.025 61.585 60.380 61.955 ;
      LAYER li1 ;
        RECT 60.660 61.945 60.830 62.135 ;
      LAYER li1 ;
        RECT 61.000 62.110 61.255 62.685 ;
      LAYER li1 ;
        RECT 60.660 61.615 60.915 61.945 ;
        RECT 46.100 61.110 46.960 61.270 ;
        RECT 45.045 60.605 45.930 60.775 ;
        RECT 46.110 60.305 46.325 60.805 ;
        RECT 46.790 60.485 46.960 61.110 ;
        RECT 47.245 60.305 47.425 61.085 ;
        RECT 48.120 60.305 48.290 61.135 ;
        RECT 48.960 60.305 49.130 61.135 ;
        RECT 49.445 60.305 54.790 61.395 ;
        RECT 54.965 60.305 58.475 61.395 ;
        RECT 59.105 60.305 59.395 61.470 ;
        RECT 60.660 61.405 60.830 61.615 ;
        RECT 60.115 61.235 60.830 61.405 ;
      LAYER li1 ;
        RECT 61.085 61.380 61.255 62.110 ;
      LAYER li1 ;
        RECT 61.430 62.015 61.690 62.855 ;
        RECT 61.865 62.085 67.210 62.855 ;
        RECT 67.385 62.105 68.595 62.855 ;
        RECT 68.855 62.305 69.025 62.595 ;
        RECT 69.195 62.475 69.525 62.855 ;
        RECT 68.855 62.135 69.520 62.305 ;
        RECT 61.865 61.565 64.445 62.085 ;
        RECT 60.115 60.475 60.285 61.235 ;
        RECT 60.500 60.305 60.830 61.065 ;
      LAYER li1 ;
        RECT 61.000 60.475 61.255 61.380 ;
      LAYER li1 ;
        RECT 61.430 60.305 61.690 61.455 ;
        RECT 64.615 61.395 67.210 61.915 ;
        RECT 67.385 61.565 67.905 62.105 ;
        RECT 68.075 61.395 68.595 61.935 ;
        RECT 61.865 60.305 67.210 61.395 ;
        RECT 67.385 60.305 68.595 61.395 ;
      LAYER li1 ;
        RECT 68.770 61.315 69.120 61.965 ;
      LAYER li1 ;
        RECT 69.290 61.145 69.520 62.135 ;
        RECT 68.855 60.975 69.520 61.145 ;
        RECT 68.855 60.475 69.025 60.975 ;
        RECT 69.195 60.305 69.525 60.805 ;
        RECT 69.695 60.475 69.920 62.595 ;
        RECT 70.135 62.395 70.385 62.855 ;
        RECT 70.570 62.405 70.900 62.575 ;
        RECT 71.080 62.405 71.830 62.575 ;
      LAYER li1 ;
        RECT 70.120 61.275 70.400 61.875 ;
      LAYER li1 ;
        RECT 70.570 60.875 70.740 62.405 ;
        RECT 70.910 61.905 71.490 62.235 ;
        RECT 70.910 61.035 71.150 61.905 ;
        RECT 71.660 61.625 71.830 62.405 ;
        RECT 72.080 62.355 72.450 62.855 ;
        RECT 72.630 62.405 73.090 62.575 ;
        RECT 73.320 62.405 73.990 62.575 ;
        RECT 72.630 62.175 72.800 62.405 ;
        RECT 72.000 61.875 72.800 62.175 ;
        RECT 72.970 61.905 73.520 62.235 ;
        RECT 72.000 61.845 72.170 61.875 ;
        RECT 72.290 61.625 72.460 61.695 ;
        RECT 71.660 61.455 72.460 61.625 ;
        RECT 71.950 61.365 72.460 61.455 ;
        RECT 71.340 60.930 71.780 61.285 ;
        RECT 70.120 60.305 70.385 60.765 ;
        RECT 70.570 60.500 70.805 60.875 ;
        RECT 71.950 60.750 72.120 61.365 ;
        RECT 71.050 60.580 72.120 60.750 ;
        RECT 72.290 60.305 72.460 61.105 ;
        RECT 72.630 60.805 72.800 61.875 ;
        RECT 72.970 60.975 73.160 61.695 ;
        RECT 73.330 61.365 73.520 61.905 ;
        RECT 73.820 61.865 73.990 62.405 ;
        RECT 74.305 62.325 74.475 62.855 ;
        RECT 74.770 62.205 75.130 62.645 ;
        RECT 75.305 62.375 75.475 62.855 ;
        RECT 76.175 62.380 76.345 62.855 ;
        RECT 77.025 62.380 77.195 62.855 ;
        RECT 74.770 62.035 75.270 62.205 ;
        RECT 75.100 61.865 75.270 62.035 ;
        RECT 77.505 62.085 82.850 62.855 ;
        RECT 83.025 62.085 86.535 62.855 ;
        RECT 87.165 62.130 87.455 62.855 ;
        RECT 87.625 62.085 92.970 62.855 ;
        RECT 93.145 62.085 98.490 62.855 ;
        RECT 98.665 62.105 99.875 62.855 ;
        RECT 73.820 61.695 74.910 61.865 ;
        RECT 75.100 61.695 76.920 61.865 ;
        RECT 73.330 61.035 73.650 61.365 ;
        RECT 72.630 60.475 72.880 60.805 ;
        RECT 73.820 60.775 73.990 61.695 ;
        RECT 75.100 61.440 75.270 61.695 ;
        RECT 77.505 61.565 80.085 62.085 ;
        RECT 74.160 61.270 75.270 61.440 ;
        RECT 80.255 61.395 82.850 61.915 ;
        RECT 83.025 61.565 84.675 62.085 ;
        RECT 84.845 61.395 86.535 61.915 ;
        RECT 87.625 61.565 90.205 62.085 ;
        RECT 74.160 61.110 75.020 61.270 ;
        RECT 73.105 60.605 73.990 60.775 ;
        RECT 74.170 60.305 74.385 60.805 ;
        RECT 74.850 60.485 75.020 61.110 ;
        RECT 75.305 60.305 75.485 61.085 ;
        RECT 76.180 60.305 76.350 61.135 ;
        RECT 77.020 60.305 77.190 61.135 ;
        RECT 77.505 60.305 82.850 61.395 ;
        RECT 83.025 60.305 86.535 61.395 ;
        RECT 87.165 60.305 87.455 61.470 ;
        RECT 90.375 61.395 92.970 61.915 ;
        RECT 93.145 61.565 95.725 62.085 ;
        RECT 95.895 61.395 98.490 61.915 ;
        RECT 87.625 60.305 92.970 61.395 ;
        RECT 93.145 60.305 98.490 61.395 ;
        RECT 98.665 61.395 99.185 61.935 ;
        RECT 99.355 61.565 99.875 62.105 ;
        RECT 98.665 60.305 99.875 61.395 ;
        RECT 16.700 60.135 16.845 60.305 ;
        RECT 17.015 60.135 17.305 60.305 ;
        RECT 17.475 60.135 17.765 60.305 ;
        RECT 17.935 60.135 18.225 60.305 ;
        RECT 18.395 60.135 18.685 60.305 ;
        RECT 18.855 60.135 19.145 60.305 ;
        RECT 19.315 60.135 19.605 60.305 ;
        RECT 19.775 60.135 20.065 60.305 ;
        RECT 20.235 60.135 20.525 60.305 ;
        RECT 20.695 60.135 20.985 60.305 ;
        RECT 21.155 60.135 21.445 60.305 ;
        RECT 21.615 60.135 21.905 60.305 ;
        RECT 22.075 60.135 22.365 60.305 ;
        RECT 22.535 60.135 22.825 60.305 ;
        RECT 22.995 60.135 23.285 60.305 ;
        RECT 23.455 60.135 23.745 60.305 ;
        RECT 23.915 60.135 24.205 60.305 ;
        RECT 24.375 60.135 24.665 60.305 ;
        RECT 24.835 60.135 25.125 60.305 ;
        RECT 25.295 60.135 25.585 60.305 ;
        RECT 25.755 60.135 26.045 60.305 ;
        RECT 26.215 60.135 26.505 60.305 ;
        RECT 26.675 60.135 26.965 60.305 ;
        RECT 27.135 60.135 27.425 60.305 ;
        RECT 27.595 60.135 27.885 60.305 ;
        RECT 28.055 60.135 28.345 60.305 ;
        RECT 28.515 60.135 28.805 60.305 ;
        RECT 28.975 60.135 29.265 60.305 ;
        RECT 29.435 60.135 29.725 60.305 ;
        RECT 29.895 60.135 30.185 60.305 ;
        RECT 30.355 60.135 30.645 60.305 ;
        RECT 30.815 60.135 31.105 60.305 ;
        RECT 31.275 60.135 31.565 60.305 ;
        RECT 31.735 60.135 32.025 60.305 ;
        RECT 32.195 60.135 32.485 60.305 ;
        RECT 32.655 60.135 32.945 60.305 ;
        RECT 33.115 60.135 33.405 60.305 ;
        RECT 33.575 60.135 33.865 60.305 ;
        RECT 34.035 60.135 34.325 60.305 ;
        RECT 34.495 60.135 34.785 60.305 ;
        RECT 34.955 60.135 35.245 60.305 ;
        RECT 35.415 60.135 35.705 60.305 ;
        RECT 35.875 60.135 36.165 60.305 ;
        RECT 36.335 60.135 36.625 60.305 ;
        RECT 36.795 60.135 37.085 60.305 ;
        RECT 37.255 60.135 37.545 60.305 ;
        RECT 37.715 60.135 38.005 60.305 ;
        RECT 38.175 60.135 38.465 60.305 ;
        RECT 38.635 60.135 38.925 60.305 ;
        RECT 39.095 60.135 39.385 60.305 ;
        RECT 39.555 60.135 39.845 60.305 ;
        RECT 40.015 60.135 40.305 60.305 ;
        RECT 40.475 60.135 40.765 60.305 ;
        RECT 40.935 60.135 41.225 60.305 ;
        RECT 41.395 60.135 41.685 60.305 ;
        RECT 41.855 60.135 42.145 60.305 ;
        RECT 42.315 60.135 42.605 60.305 ;
        RECT 42.775 60.135 43.065 60.305 ;
        RECT 43.235 60.135 43.525 60.305 ;
        RECT 43.695 60.135 43.985 60.305 ;
        RECT 44.155 60.135 44.445 60.305 ;
        RECT 44.615 60.135 44.905 60.305 ;
        RECT 45.075 60.135 45.365 60.305 ;
        RECT 45.535 60.135 45.825 60.305 ;
        RECT 45.995 60.135 46.285 60.305 ;
        RECT 46.455 60.135 46.745 60.305 ;
        RECT 46.915 60.135 47.205 60.305 ;
        RECT 47.375 60.135 47.665 60.305 ;
        RECT 47.835 60.135 48.125 60.305 ;
        RECT 48.295 60.135 48.585 60.305 ;
        RECT 48.755 60.135 49.045 60.305 ;
        RECT 49.215 60.135 49.505 60.305 ;
        RECT 49.675 60.135 49.965 60.305 ;
        RECT 50.135 60.135 50.425 60.305 ;
        RECT 50.595 60.135 50.885 60.305 ;
        RECT 51.055 60.135 51.345 60.305 ;
        RECT 51.515 60.135 51.805 60.305 ;
        RECT 51.975 60.135 52.265 60.305 ;
        RECT 52.435 60.135 52.725 60.305 ;
        RECT 52.895 60.135 53.185 60.305 ;
        RECT 53.355 60.135 53.645 60.305 ;
        RECT 53.815 60.135 54.105 60.305 ;
        RECT 54.275 60.135 54.565 60.305 ;
        RECT 54.735 60.135 55.025 60.305 ;
        RECT 55.195 60.135 55.485 60.305 ;
        RECT 55.655 60.135 55.945 60.305 ;
        RECT 56.115 60.135 56.405 60.305 ;
        RECT 56.575 60.135 56.865 60.305 ;
        RECT 57.035 60.135 57.325 60.305 ;
        RECT 57.495 60.135 57.785 60.305 ;
        RECT 57.955 60.135 58.245 60.305 ;
        RECT 58.415 60.135 58.705 60.305 ;
        RECT 58.875 60.135 59.165 60.305 ;
        RECT 59.335 60.135 59.625 60.305 ;
        RECT 59.795 60.135 60.085 60.305 ;
        RECT 60.255 60.135 60.545 60.305 ;
        RECT 60.715 60.135 61.005 60.305 ;
        RECT 61.175 60.135 61.465 60.305 ;
        RECT 61.635 60.135 61.925 60.305 ;
        RECT 62.095 60.135 62.385 60.305 ;
        RECT 62.555 60.135 62.845 60.305 ;
        RECT 63.015 60.135 63.305 60.305 ;
        RECT 63.475 60.135 63.765 60.305 ;
        RECT 63.935 60.135 64.225 60.305 ;
        RECT 64.395 60.135 64.685 60.305 ;
        RECT 64.855 60.135 65.145 60.305 ;
        RECT 65.315 60.135 65.605 60.305 ;
        RECT 65.775 60.135 66.065 60.305 ;
        RECT 66.235 60.135 66.525 60.305 ;
        RECT 66.695 60.135 66.985 60.305 ;
        RECT 67.155 60.135 67.445 60.305 ;
        RECT 67.615 60.135 67.905 60.305 ;
        RECT 68.075 60.135 68.365 60.305 ;
        RECT 68.535 60.135 68.825 60.305 ;
        RECT 68.995 60.135 69.285 60.305 ;
        RECT 69.455 60.135 69.745 60.305 ;
        RECT 69.915 60.135 70.205 60.305 ;
        RECT 70.375 60.135 70.665 60.305 ;
        RECT 70.835 60.135 71.125 60.305 ;
        RECT 71.295 60.135 71.585 60.305 ;
        RECT 71.755 60.135 72.045 60.305 ;
        RECT 72.215 60.135 72.505 60.305 ;
        RECT 72.675 60.135 72.965 60.305 ;
        RECT 73.135 60.135 73.425 60.305 ;
        RECT 73.595 60.135 73.885 60.305 ;
        RECT 74.055 60.135 74.345 60.305 ;
        RECT 74.515 60.135 74.805 60.305 ;
        RECT 74.975 60.135 75.265 60.305 ;
        RECT 75.435 60.135 75.725 60.305 ;
        RECT 75.895 60.135 76.185 60.305 ;
        RECT 76.355 60.135 76.645 60.305 ;
        RECT 76.815 60.135 77.105 60.305 ;
        RECT 77.275 60.135 77.565 60.305 ;
        RECT 77.735 60.135 78.025 60.305 ;
        RECT 78.195 60.135 78.485 60.305 ;
        RECT 78.655 60.135 78.945 60.305 ;
        RECT 79.115 60.135 79.405 60.305 ;
        RECT 79.575 60.135 79.865 60.305 ;
        RECT 80.035 60.135 80.325 60.305 ;
        RECT 80.495 60.135 80.785 60.305 ;
        RECT 80.955 60.135 81.245 60.305 ;
        RECT 81.415 60.135 81.705 60.305 ;
        RECT 81.875 60.135 82.165 60.305 ;
        RECT 82.335 60.135 82.625 60.305 ;
        RECT 82.795 60.135 83.085 60.305 ;
        RECT 83.255 60.135 83.545 60.305 ;
        RECT 83.715 60.135 84.005 60.305 ;
        RECT 84.175 60.135 84.465 60.305 ;
        RECT 84.635 60.135 84.925 60.305 ;
        RECT 85.095 60.135 85.385 60.305 ;
        RECT 85.555 60.135 85.845 60.305 ;
        RECT 86.015 60.135 86.305 60.305 ;
        RECT 86.475 60.135 86.765 60.305 ;
        RECT 86.935 60.135 87.225 60.305 ;
        RECT 87.395 60.135 87.685 60.305 ;
        RECT 87.855 60.135 88.145 60.305 ;
        RECT 88.315 60.135 88.605 60.305 ;
        RECT 88.775 60.135 89.065 60.305 ;
        RECT 89.235 60.135 89.525 60.305 ;
        RECT 89.695 60.135 89.985 60.305 ;
        RECT 90.155 60.135 90.445 60.305 ;
        RECT 90.615 60.135 90.905 60.305 ;
        RECT 91.075 60.135 91.365 60.305 ;
        RECT 91.535 60.135 91.825 60.305 ;
        RECT 91.995 60.135 92.285 60.305 ;
        RECT 92.455 60.135 92.745 60.305 ;
        RECT 92.915 60.135 93.205 60.305 ;
        RECT 93.375 60.135 93.665 60.305 ;
        RECT 93.835 60.135 94.125 60.305 ;
        RECT 94.295 60.135 94.585 60.305 ;
        RECT 94.755 60.135 95.045 60.305 ;
        RECT 95.215 60.135 95.505 60.305 ;
        RECT 95.675 60.135 95.965 60.305 ;
        RECT 96.135 60.135 96.425 60.305 ;
        RECT 96.595 60.135 96.885 60.305 ;
        RECT 97.055 60.135 97.345 60.305 ;
        RECT 97.515 60.135 97.805 60.305 ;
        RECT 97.975 60.135 98.265 60.305 ;
        RECT 98.435 60.135 98.725 60.305 ;
        RECT 98.895 60.135 99.185 60.305 ;
        RECT 99.355 60.135 99.645 60.305 ;
        RECT 99.815 60.135 99.960 60.305 ;
        RECT 16.785 59.045 17.995 60.135 ;
        RECT 18.165 59.045 23.510 60.135 ;
        RECT 23.685 59.045 29.030 60.135 ;
        RECT 29.205 59.045 34.550 60.135 ;
        RECT 34.725 59.045 37.315 60.135 ;
        RECT 37.955 59.380 38.285 60.135 ;
        RECT 38.465 59.250 38.645 59.965 ;
        RECT 38.850 59.435 39.180 60.135 ;
      LAYER li1 ;
        RECT 39.390 59.260 39.580 59.965 ;
      LAYER li1 ;
        RECT 39.750 59.435 40.080 60.135 ;
      LAYER li1 ;
        RECT 40.250 59.265 40.440 59.965 ;
      LAYER li1 ;
        RECT 40.610 59.435 40.940 60.135 ;
      LAYER li1 ;
        RECT 40.250 59.260 40.995 59.265 ;
      LAYER li1 ;
        RECT 38.465 59.080 39.220 59.250 ;
        RECT 16.785 58.335 17.305 58.875 ;
        RECT 17.475 58.505 17.995 59.045 ;
        RECT 18.165 58.355 20.745 58.875 ;
        RECT 20.915 58.525 23.510 59.045 ;
        RECT 23.685 58.355 26.265 58.875 ;
        RECT 26.435 58.525 29.030 59.045 ;
        RECT 29.205 58.355 31.785 58.875 ;
        RECT 31.955 58.525 34.550 59.045 ;
        RECT 34.725 58.355 35.935 58.875 ;
        RECT 36.105 58.525 37.315 59.045 ;
        RECT 39.010 58.855 39.220 59.080 ;
      LAYER li1 ;
        RECT 39.390 59.035 40.995 59.260 ;
      LAYER li1 ;
        RECT 41.165 59.045 44.675 60.135 ;
      LAYER li1 ;
        RECT 38.465 58.495 38.840 58.825 ;
      LAYER li1 ;
        RECT 39.010 58.520 40.545 58.855 ;
        RECT 16.785 57.585 17.995 58.335 ;
        RECT 18.165 57.585 23.510 58.355 ;
        RECT 23.685 57.585 29.030 58.355 ;
        RECT 29.205 57.585 34.550 58.355 ;
        RECT 34.725 57.585 37.315 58.355 ;
        RECT 39.010 58.305 39.220 58.520 ;
      LAYER li1 ;
        RECT 40.715 58.345 40.995 59.035 ;
      LAYER li1 ;
        RECT 37.955 58.115 39.220 58.305 ;
      LAYER li1 ;
        RECT 39.390 58.115 40.995 58.345 ;
      LAYER li1 ;
        RECT 41.165 58.355 42.815 58.875 ;
        RECT 42.985 58.525 44.675 59.045 ;
        RECT 44.845 58.970 45.135 60.135 ;
        RECT 45.305 59.045 50.650 60.135 ;
        RECT 50.825 59.045 56.170 60.135 ;
        RECT 56.345 59.045 61.690 60.135 ;
        RECT 61.865 59.045 63.535 60.135 ;
        RECT 63.715 59.380 64.045 60.135 ;
        RECT 64.225 59.250 64.405 59.965 ;
        RECT 64.610 59.435 64.940 60.135 ;
      LAYER li1 ;
        RECT 65.150 59.795 65.340 59.965 ;
        RECT 65.145 59.625 65.340 59.795 ;
        RECT 65.150 59.260 65.340 59.625 ;
      LAYER li1 ;
        RECT 65.510 59.435 65.840 60.135 ;
      LAYER li1 ;
        RECT 66.010 59.265 66.200 59.965 ;
      LAYER li1 ;
        RECT 66.370 59.435 66.700 60.135 ;
      LAYER li1 ;
        RECT 66.010 59.260 66.755 59.265 ;
      LAYER li1 ;
        RECT 45.305 58.355 47.885 58.875 ;
        RECT 48.055 58.525 50.650 59.045 ;
        RECT 50.825 58.355 53.405 58.875 ;
        RECT 53.575 58.525 56.170 59.045 ;
        RECT 56.345 58.355 58.925 58.875 ;
        RECT 59.095 58.525 61.690 59.045 ;
        RECT 61.865 58.355 62.615 58.875 ;
        RECT 62.785 58.525 63.535 59.045 ;
      LAYER li1 ;
        RECT 63.745 58.495 64.055 59.115 ;
      LAYER li1 ;
        RECT 64.225 59.080 64.980 59.250 ;
        RECT 64.770 58.855 64.980 59.080 ;
      LAYER li1 ;
        RECT 65.150 59.035 66.755 59.260 ;
      LAYER li1 ;
        RECT 66.925 59.045 72.270 60.135 ;
        RECT 64.770 58.520 66.305 58.855 ;
        RECT 37.955 57.755 38.285 58.115 ;
      LAYER li1 ;
        RECT 39.390 58.015 39.580 58.115 ;
      LAYER li1 ;
        RECT 38.815 57.585 39.145 57.945 ;
        RECT 39.750 57.585 40.080 57.945 ;
      LAYER li1 ;
        RECT 40.250 57.755 40.440 58.115 ;
      LAYER li1 ;
        RECT 40.610 57.585 40.940 57.945 ;
        RECT 41.165 57.585 44.675 58.355 ;
        RECT 44.845 57.585 45.135 58.310 ;
        RECT 45.305 57.585 50.650 58.355 ;
        RECT 50.825 57.585 56.170 58.355 ;
        RECT 56.345 57.585 61.690 58.355 ;
        RECT 61.865 57.585 63.535 58.355 ;
        RECT 64.770 58.305 64.980 58.520 ;
      LAYER li1 ;
        RECT 66.475 58.345 66.755 59.035 ;
      LAYER li1 ;
        RECT 63.715 58.115 64.980 58.305 ;
      LAYER li1 ;
        RECT 65.150 58.115 66.755 58.345 ;
      LAYER li1 ;
        RECT 66.925 58.355 69.505 58.875 ;
        RECT 69.675 58.525 72.270 59.045 ;
        RECT 72.905 58.970 73.195 60.135 ;
        RECT 73.365 59.045 78.710 60.135 ;
        RECT 78.885 59.045 84.230 60.135 ;
        RECT 84.405 59.045 89.750 60.135 ;
        RECT 89.925 59.045 95.270 60.135 ;
        RECT 95.445 59.045 98.035 60.135 ;
        RECT 73.365 58.355 75.945 58.875 ;
        RECT 76.115 58.525 78.710 59.045 ;
        RECT 78.885 58.355 81.465 58.875 ;
        RECT 81.635 58.525 84.230 59.045 ;
        RECT 84.405 58.355 86.985 58.875 ;
        RECT 87.155 58.525 89.750 59.045 ;
        RECT 89.925 58.355 92.505 58.875 ;
        RECT 92.675 58.525 95.270 59.045 ;
        RECT 95.445 58.355 96.655 58.875 ;
        RECT 96.825 58.525 98.035 59.045 ;
        RECT 98.665 59.045 99.875 60.135 ;
        RECT 98.665 58.505 99.185 59.045 ;
        RECT 63.715 57.755 64.045 58.115 ;
      LAYER li1 ;
        RECT 65.150 58.015 65.340 58.115 ;
      LAYER li1 ;
        RECT 64.575 57.585 64.905 57.945 ;
        RECT 65.510 57.585 65.840 57.945 ;
      LAYER li1 ;
        RECT 66.010 57.755 66.200 58.115 ;
      LAYER li1 ;
        RECT 66.370 57.585 66.700 57.945 ;
        RECT 66.925 57.585 72.270 58.355 ;
        RECT 72.905 57.585 73.195 58.310 ;
        RECT 73.365 57.585 78.710 58.355 ;
        RECT 78.885 57.585 84.230 58.355 ;
        RECT 84.405 57.585 89.750 58.355 ;
        RECT 89.925 57.585 95.270 58.355 ;
        RECT 95.445 57.585 98.035 58.355 ;
        RECT 99.355 58.335 99.875 58.875 ;
        RECT 98.665 57.585 99.875 58.335 ;
        RECT 16.700 57.415 16.845 57.585 ;
        RECT 17.015 57.415 17.305 57.585 ;
        RECT 17.475 57.415 17.765 57.585 ;
        RECT 17.935 57.415 18.225 57.585 ;
        RECT 18.395 57.415 18.685 57.585 ;
        RECT 18.855 57.415 19.145 57.585 ;
        RECT 19.315 57.415 19.605 57.585 ;
        RECT 19.775 57.415 20.065 57.585 ;
        RECT 20.235 57.415 20.525 57.585 ;
        RECT 20.695 57.415 20.985 57.585 ;
        RECT 21.155 57.415 21.445 57.585 ;
        RECT 21.615 57.415 21.905 57.585 ;
        RECT 22.075 57.415 22.365 57.585 ;
        RECT 22.535 57.415 22.825 57.585 ;
        RECT 22.995 57.415 23.285 57.585 ;
        RECT 23.455 57.415 23.745 57.585 ;
        RECT 23.915 57.415 24.205 57.585 ;
        RECT 24.375 57.415 24.665 57.585 ;
        RECT 24.835 57.415 25.125 57.585 ;
        RECT 25.295 57.415 25.585 57.585 ;
        RECT 25.755 57.415 26.045 57.585 ;
        RECT 26.215 57.415 26.505 57.585 ;
        RECT 26.675 57.415 26.965 57.585 ;
        RECT 27.135 57.415 27.425 57.585 ;
        RECT 27.595 57.415 27.885 57.585 ;
        RECT 28.055 57.415 28.345 57.585 ;
        RECT 28.515 57.415 28.805 57.585 ;
        RECT 28.975 57.415 29.265 57.585 ;
        RECT 29.435 57.415 29.725 57.585 ;
        RECT 29.895 57.415 30.185 57.585 ;
        RECT 30.355 57.415 30.645 57.585 ;
        RECT 30.815 57.415 31.105 57.585 ;
        RECT 31.275 57.415 31.565 57.585 ;
        RECT 31.735 57.415 32.025 57.585 ;
        RECT 32.195 57.415 32.485 57.585 ;
        RECT 32.655 57.415 32.945 57.585 ;
        RECT 33.115 57.415 33.405 57.585 ;
        RECT 33.575 57.415 33.865 57.585 ;
        RECT 34.035 57.415 34.325 57.585 ;
        RECT 34.495 57.415 34.785 57.585 ;
        RECT 34.955 57.415 35.245 57.585 ;
        RECT 35.415 57.415 35.705 57.585 ;
        RECT 35.875 57.415 36.165 57.585 ;
        RECT 36.335 57.415 36.625 57.585 ;
        RECT 36.795 57.415 37.085 57.585 ;
        RECT 37.255 57.415 37.545 57.585 ;
        RECT 37.715 57.415 38.005 57.585 ;
        RECT 38.175 57.415 38.465 57.585 ;
        RECT 38.635 57.415 38.925 57.585 ;
        RECT 39.095 57.415 39.385 57.585 ;
        RECT 39.555 57.415 39.845 57.585 ;
        RECT 40.015 57.415 40.305 57.585 ;
        RECT 40.475 57.415 40.765 57.585 ;
        RECT 40.935 57.415 41.225 57.585 ;
        RECT 41.395 57.415 41.685 57.585 ;
        RECT 41.855 57.415 42.145 57.585 ;
        RECT 42.315 57.415 42.605 57.585 ;
        RECT 42.775 57.415 43.065 57.585 ;
        RECT 43.235 57.415 43.525 57.585 ;
        RECT 43.695 57.415 43.985 57.585 ;
        RECT 44.155 57.415 44.445 57.585 ;
        RECT 44.615 57.415 44.905 57.585 ;
        RECT 45.075 57.415 45.365 57.585 ;
        RECT 45.535 57.415 45.825 57.585 ;
        RECT 45.995 57.415 46.285 57.585 ;
        RECT 46.455 57.415 46.745 57.585 ;
        RECT 46.915 57.415 47.205 57.585 ;
        RECT 47.375 57.415 47.665 57.585 ;
        RECT 47.835 57.415 48.125 57.585 ;
        RECT 48.295 57.415 48.585 57.585 ;
        RECT 48.755 57.415 49.045 57.585 ;
        RECT 49.215 57.415 49.505 57.585 ;
        RECT 49.675 57.415 49.965 57.585 ;
        RECT 50.135 57.415 50.425 57.585 ;
        RECT 50.595 57.415 50.885 57.585 ;
        RECT 51.055 57.415 51.345 57.585 ;
        RECT 51.515 57.415 51.805 57.585 ;
        RECT 51.975 57.415 52.265 57.585 ;
        RECT 52.435 57.415 52.725 57.585 ;
        RECT 52.895 57.415 53.185 57.585 ;
        RECT 53.355 57.415 53.645 57.585 ;
        RECT 53.815 57.415 54.105 57.585 ;
        RECT 54.275 57.415 54.565 57.585 ;
        RECT 54.735 57.415 55.025 57.585 ;
        RECT 55.195 57.415 55.485 57.585 ;
        RECT 55.655 57.415 55.945 57.585 ;
        RECT 56.115 57.415 56.405 57.585 ;
        RECT 56.575 57.415 56.865 57.585 ;
        RECT 57.035 57.415 57.325 57.585 ;
        RECT 57.495 57.415 57.785 57.585 ;
        RECT 57.955 57.415 58.245 57.585 ;
        RECT 58.415 57.415 58.705 57.585 ;
        RECT 58.875 57.415 59.165 57.585 ;
        RECT 59.335 57.415 59.625 57.585 ;
        RECT 59.795 57.415 60.085 57.585 ;
        RECT 60.255 57.415 60.545 57.585 ;
        RECT 60.715 57.415 61.005 57.585 ;
        RECT 61.175 57.415 61.465 57.585 ;
        RECT 61.635 57.415 61.925 57.585 ;
        RECT 62.095 57.415 62.385 57.585 ;
        RECT 62.555 57.415 62.845 57.585 ;
        RECT 63.015 57.415 63.305 57.585 ;
        RECT 63.475 57.415 63.765 57.585 ;
        RECT 63.935 57.415 64.225 57.585 ;
        RECT 64.395 57.415 64.685 57.585 ;
        RECT 64.855 57.415 65.145 57.585 ;
        RECT 65.315 57.415 65.605 57.585 ;
        RECT 65.775 57.415 66.065 57.585 ;
        RECT 66.235 57.415 66.525 57.585 ;
        RECT 66.695 57.415 66.985 57.585 ;
        RECT 67.155 57.415 67.445 57.585 ;
        RECT 67.615 57.415 67.905 57.585 ;
        RECT 68.075 57.415 68.365 57.585 ;
        RECT 68.535 57.415 68.825 57.585 ;
        RECT 68.995 57.415 69.285 57.585 ;
        RECT 69.455 57.415 69.745 57.585 ;
        RECT 69.915 57.415 70.205 57.585 ;
        RECT 70.375 57.415 70.665 57.585 ;
        RECT 70.835 57.415 71.125 57.585 ;
        RECT 71.295 57.415 71.585 57.585 ;
        RECT 71.755 57.415 72.045 57.585 ;
        RECT 72.215 57.415 72.505 57.585 ;
        RECT 72.675 57.415 72.965 57.585 ;
        RECT 73.135 57.415 73.425 57.585 ;
        RECT 73.595 57.415 73.885 57.585 ;
        RECT 74.055 57.415 74.345 57.585 ;
        RECT 74.515 57.415 74.805 57.585 ;
        RECT 74.975 57.415 75.265 57.585 ;
        RECT 75.435 57.415 75.725 57.585 ;
        RECT 75.895 57.415 76.185 57.585 ;
        RECT 76.355 57.415 76.645 57.585 ;
        RECT 76.815 57.415 77.105 57.585 ;
        RECT 77.275 57.415 77.565 57.585 ;
        RECT 77.735 57.415 78.025 57.585 ;
        RECT 78.195 57.415 78.485 57.585 ;
        RECT 78.655 57.415 78.945 57.585 ;
        RECT 79.115 57.415 79.405 57.585 ;
        RECT 79.575 57.415 79.865 57.585 ;
        RECT 80.035 57.415 80.325 57.585 ;
        RECT 80.495 57.415 80.785 57.585 ;
        RECT 80.955 57.415 81.245 57.585 ;
        RECT 81.415 57.415 81.705 57.585 ;
        RECT 81.875 57.415 82.165 57.585 ;
        RECT 82.335 57.415 82.625 57.585 ;
        RECT 82.795 57.415 83.085 57.585 ;
        RECT 83.255 57.415 83.545 57.585 ;
        RECT 83.715 57.415 84.005 57.585 ;
        RECT 84.175 57.415 84.465 57.585 ;
        RECT 84.635 57.415 84.925 57.585 ;
        RECT 85.095 57.415 85.385 57.585 ;
        RECT 85.555 57.415 85.845 57.585 ;
        RECT 86.015 57.415 86.305 57.585 ;
        RECT 86.475 57.415 86.765 57.585 ;
        RECT 86.935 57.415 87.225 57.585 ;
        RECT 87.395 57.415 87.685 57.585 ;
        RECT 87.855 57.415 88.145 57.585 ;
        RECT 88.315 57.415 88.605 57.585 ;
        RECT 88.775 57.415 89.065 57.585 ;
        RECT 89.235 57.415 89.525 57.585 ;
        RECT 89.695 57.415 89.985 57.585 ;
        RECT 90.155 57.415 90.445 57.585 ;
        RECT 90.615 57.415 90.905 57.585 ;
        RECT 91.075 57.415 91.365 57.585 ;
        RECT 91.535 57.415 91.825 57.585 ;
        RECT 91.995 57.415 92.285 57.585 ;
        RECT 92.455 57.415 92.745 57.585 ;
        RECT 92.915 57.415 93.205 57.585 ;
        RECT 93.375 57.415 93.665 57.585 ;
        RECT 93.835 57.415 94.125 57.585 ;
        RECT 94.295 57.415 94.585 57.585 ;
        RECT 94.755 57.415 95.045 57.585 ;
        RECT 95.215 57.415 95.505 57.585 ;
        RECT 95.675 57.415 95.965 57.585 ;
        RECT 96.135 57.415 96.425 57.585 ;
        RECT 96.595 57.415 96.885 57.585 ;
        RECT 97.055 57.415 97.345 57.585 ;
        RECT 97.515 57.415 97.805 57.585 ;
        RECT 97.975 57.415 98.265 57.585 ;
        RECT 98.435 57.415 98.725 57.585 ;
        RECT 98.895 57.415 99.185 57.585 ;
        RECT 99.355 57.415 99.645 57.585 ;
        RECT 99.815 57.415 99.960 57.585 ;
        RECT 16.785 56.665 17.995 57.415 ;
        RECT 16.785 56.125 17.305 56.665 ;
        RECT 18.165 56.645 23.510 57.415 ;
        RECT 23.685 56.645 29.030 57.415 ;
        RECT 29.205 56.645 30.875 57.415 ;
        RECT 31.045 56.690 31.335 57.415 ;
        RECT 31.505 56.645 36.850 57.415 ;
        RECT 37.025 56.645 42.370 57.415 ;
        RECT 42.545 56.645 47.890 57.415 ;
        RECT 48.065 56.645 53.410 57.415 ;
        RECT 53.585 56.645 58.930 57.415 ;
        RECT 59.105 56.690 59.395 57.415 ;
        RECT 59.565 56.645 64.910 57.415 ;
        RECT 65.095 56.885 65.425 57.245 ;
        RECT 65.955 57.055 66.285 57.415 ;
        RECT 66.890 57.055 67.220 57.415 ;
      LAYER li1 ;
        RECT 66.530 56.885 66.720 56.985 ;
        RECT 67.390 56.885 67.580 57.245 ;
      LAYER li1 ;
        RECT 67.750 57.055 68.080 57.415 ;
        RECT 65.095 56.695 66.360 56.885 ;
        RECT 17.475 55.955 17.995 56.495 ;
        RECT 18.165 56.125 20.745 56.645 ;
        RECT 20.915 55.955 23.510 56.475 ;
        RECT 23.685 56.125 26.265 56.645 ;
        RECT 26.435 55.955 29.030 56.475 ;
        RECT 29.205 56.125 29.955 56.645 ;
        RECT 30.125 55.955 30.875 56.475 ;
        RECT 31.505 56.125 34.085 56.645 ;
        RECT 16.785 54.865 17.995 55.955 ;
        RECT 18.165 54.865 23.510 55.955 ;
        RECT 23.685 54.865 29.030 55.955 ;
        RECT 29.205 54.865 30.875 55.955 ;
        RECT 31.045 54.865 31.335 56.030 ;
        RECT 34.255 55.955 36.850 56.475 ;
        RECT 37.025 56.125 39.605 56.645 ;
        RECT 39.775 55.955 42.370 56.475 ;
        RECT 42.545 56.125 45.125 56.645 ;
        RECT 45.295 55.955 47.890 56.475 ;
        RECT 48.065 56.125 50.645 56.645 ;
        RECT 50.815 55.955 53.410 56.475 ;
        RECT 53.585 56.125 56.165 56.645 ;
        RECT 56.335 55.955 58.930 56.475 ;
        RECT 59.565 56.125 62.145 56.645 ;
        RECT 31.505 54.865 36.850 55.955 ;
        RECT 37.025 54.865 42.370 55.955 ;
        RECT 42.545 54.865 47.890 55.955 ;
        RECT 48.065 54.865 53.410 55.955 ;
        RECT 53.585 54.865 58.930 55.955 ;
        RECT 59.105 54.865 59.395 56.030 ;
        RECT 62.315 55.955 64.910 56.475 ;
        RECT 59.565 54.865 64.910 55.955 ;
      LAYER li1 ;
        RECT 65.125 55.885 65.435 56.505 ;
      LAYER li1 ;
        RECT 66.150 56.480 66.360 56.695 ;
      LAYER li1 ;
        RECT 66.530 56.655 68.135 56.885 ;
      LAYER li1 ;
        RECT 66.150 56.145 67.685 56.480 ;
        RECT 66.150 55.920 66.360 56.145 ;
      LAYER li1 ;
        RECT 67.855 55.965 68.135 56.655 ;
      LAYER li1 ;
        RECT 68.305 56.645 73.650 57.415 ;
        RECT 73.825 56.645 79.170 57.415 ;
        RECT 79.345 56.645 84.690 57.415 ;
        RECT 84.865 56.645 86.535 57.415 ;
        RECT 87.165 56.690 87.455 57.415 ;
        RECT 87.625 56.645 92.970 57.415 ;
        RECT 93.145 56.645 98.490 57.415 ;
        RECT 98.665 56.665 99.875 57.415 ;
        RECT 68.305 56.125 70.885 56.645 ;
        RECT 65.605 55.750 66.360 55.920 ;
        RECT 65.095 54.865 65.425 55.620 ;
        RECT 65.605 55.035 65.785 55.750 ;
      LAYER li1 ;
        RECT 66.530 55.740 68.135 55.965 ;
      LAYER li1 ;
        RECT 71.055 55.955 73.650 56.475 ;
        RECT 73.825 56.125 76.405 56.645 ;
        RECT 76.575 55.955 79.170 56.475 ;
        RECT 79.345 56.125 81.925 56.645 ;
        RECT 82.095 55.955 84.690 56.475 ;
        RECT 84.865 56.125 85.615 56.645 ;
        RECT 85.785 55.955 86.535 56.475 ;
        RECT 87.625 56.125 90.205 56.645 ;
        RECT 65.990 54.865 66.320 55.565 ;
      LAYER li1 ;
        RECT 66.530 55.035 66.720 55.740 ;
        RECT 67.390 55.735 68.135 55.740 ;
      LAYER li1 ;
        RECT 66.890 54.865 67.220 55.565 ;
      LAYER li1 ;
        RECT 67.390 55.035 67.580 55.735 ;
      LAYER li1 ;
        RECT 67.750 54.865 68.080 55.565 ;
        RECT 68.305 54.865 73.650 55.955 ;
        RECT 73.825 54.865 79.170 55.955 ;
        RECT 79.345 54.865 84.690 55.955 ;
        RECT 84.865 54.865 86.535 55.955 ;
        RECT 87.165 54.865 87.455 56.030 ;
        RECT 90.375 55.955 92.970 56.475 ;
        RECT 93.145 56.125 95.725 56.645 ;
        RECT 95.895 55.955 98.490 56.475 ;
        RECT 87.625 54.865 92.970 55.955 ;
        RECT 93.145 54.865 98.490 55.955 ;
        RECT 98.665 55.955 99.185 56.495 ;
        RECT 99.355 56.125 99.875 56.665 ;
        RECT 98.665 54.865 99.875 55.955 ;
        RECT 16.700 54.695 16.845 54.865 ;
        RECT 17.015 54.695 17.305 54.865 ;
        RECT 17.475 54.695 17.765 54.865 ;
        RECT 17.935 54.695 18.225 54.865 ;
        RECT 18.395 54.695 18.685 54.865 ;
        RECT 18.855 54.695 19.145 54.865 ;
        RECT 19.315 54.695 19.605 54.865 ;
        RECT 19.775 54.695 20.065 54.865 ;
        RECT 20.235 54.695 20.525 54.865 ;
        RECT 20.695 54.695 20.985 54.865 ;
        RECT 21.155 54.695 21.445 54.865 ;
        RECT 21.615 54.695 21.905 54.865 ;
        RECT 22.075 54.695 22.365 54.865 ;
        RECT 22.535 54.695 22.825 54.865 ;
        RECT 22.995 54.695 23.285 54.865 ;
        RECT 23.455 54.695 23.745 54.865 ;
        RECT 23.915 54.695 24.205 54.865 ;
        RECT 24.375 54.695 24.665 54.865 ;
        RECT 24.835 54.695 25.125 54.865 ;
        RECT 25.295 54.695 25.585 54.865 ;
        RECT 25.755 54.695 26.045 54.865 ;
        RECT 26.215 54.695 26.505 54.865 ;
        RECT 26.675 54.695 26.965 54.865 ;
        RECT 27.135 54.695 27.425 54.865 ;
        RECT 27.595 54.695 27.885 54.865 ;
        RECT 28.055 54.695 28.345 54.865 ;
        RECT 28.515 54.695 28.805 54.865 ;
        RECT 28.975 54.695 29.265 54.865 ;
        RECT 29.435 54.695 29.725 54.865 ;
        RECT 29.895 54.695 30.185 54.865 ;
        RECT 30.355 54.695 30.645 54.865 ;
        RECT 30.815 54.695 31.105 54.865 ;
        RECT 31.275 54.695 31.565 54.865 ;
        RECT 31.735 54.695 32.025 54.865 ;
        RECT 32.195 54.695 32.485 54.865 ;
        RECT 32.655 54.695 32.945 54.865 ;
        RECT 33.115 54.695 33.405 54.865 ;
        RECT 33.575 54.695 33.865 54.865 ;
        RECT 34.035 54.695 34.325 54.865 ;
        RECT 34.495 54.695 34.785 54.865 ;
        RECT 34.955 54.695 35.245 54.865 ;
        RECT 35.415 54.695 35.705 54.865 ;
        RECT 35.875 54.695 36.165 54.865 ;
        RECT 36.335 54.695 36.625 54.865 ;
        RECT 36.795 54.695 37.085 54.865 ;
        RECT 37.255 54.695 37.545 54.865 ;
        RECT 37.715 54.695 38.005 54.865 ;
        RECT 38.175 54.695 38.465 54.865 ;
        RECT 38.635 54.695 38.925 54.865 ;
        RECT 39.095 54.695 39.385 54.865 ;
        RECT 39.555 54.695 39.845 54.865 ;
        RECT 40.015 54.695 40.305 54.865 ;
        RECT 40.475 54.695 40.765 54.865 ;
        RECT 40.935 54.695 41.225 54.865 ;
        RECT 41.395 54.695 41.685 54.865 ;
        RECT 41.855 54.695 42.145 54.865 ;
        RECT 42.315 54.695 42.605 54.865 ;
        RECT 42.775 54.695 43.065 54.865 ;
        RECT 43.235 54.695 43.525 54.865 ;
        RECT 43.695 54.695 43.985 54.865 ;
        RECT 44.155 54.695 44.445 54.865 ;
        RECT 44.615 54.695 44.905 54.865 ;
        RECT 45.075 54.695 45.365 54.865 ;
        RECT 45.535 54.695 45.825 54.865 ;
        RECT 45.995 54.695 46.285 54.865 ;
        RECT 46.455 54.695 46.745 54.865 ;
        RECT 46.915 54.695 47.205 54.865 ;
        RECT 47.375 54.695 47.665 54.865 ;
        RECT 47.835 54.695 48.125 54.865 ;
        RECT 48.295 54.695 48.585 54.865 ;
        RECT 48.755 54.695 49.045 54.865 ;
        RECT 49.215 54.695 49.505 54.865 ;
        RECT 49.675 54.695 49.965 54.865 ;
        RECT 50.135 54.695 50.425 54.865 ;
        RECT 50.595 54.695 50.885 54.865 ;
        RECT 51.055 54.695 51.345 54.865 ;
        RECT 51.515 54.695 51.805 54.865 ;
        RECT 51.975 54.695 52.265 54.865 ;
        RECT 52.435 54.695 52.725 54.865 ;
        RECT 52.895 54.695 53.185 54.865 ;
        RECT 53.355 54.695 53.645 54.865 ;
        RECT 53.815 54.695 54.105 54.865 ;
        RECT 54.275 54.695 54.565 54.865 ;
        RECT 54.735 54.695 55.025 54.865 ;
        RECT 55.195 54.695 55.485 54.865 ;
        RECT 55.655 54.695 55.945 54.865 ;
        RECT 56.115 54.695 56.405 54.865 ;
        RECT 56.575 54.695 56.865 54.865 ;
        RECT 57.035 54.695 57.325 54.865 ;
        RECT 57.495 54.695 57.785 54.865 ;
        RECT 57.955 54.695 58.245 54.865 ;
        RECT 58.415 54.695 58.705 54.865 ;
        RECT 58.875 54.695 59.165 54.865 ;
        RECT 59.335 54.695 59.625 54.865 ;
        RECT 59.795 54.695 60.085 54.865 ;
        RECT 60.255 54.695 60.545 54.865 ;
        RECT 60.715 54.695 61.005 54.865 ;
        RECT 61.175 54.695 61.465 54.865 ;
        RECT 61.635 54.695 61.925 54.865 ;
        RECT 62.095 54.695 62.385 54.865 ;
        RECT 62.555 54.695 62.845 54.865 ;
        RECT 63.015 54.695 63.305 54.865 ;
        RECT 63.475 54.695 63.765 54.865 ;
        RECT 63.935 54.695 64.225 54.865 ;
        RECT 64.395 54.695 64.685 54.865 ;
        RECT 64.855 54.695 65.145 54.865 ;
        RECT 65.315 54.695 65.605 54.865 ;
        RECT 65.775 54.695 66.065 54.865 ;
        RECT 66.235 54.695 66.525 54.865 ;
        RECT 66.695 54.695 66.985 54.865 ;
        RECT 67.155 54.695 67.445 54.865 ;
        RECT 67.615 54.695 67.905 54.865 ;
        RECT 68.075 54.695 68.365 54.865 ;
        RECT 68.535 54.695 68.825 54.865 ;
        RECT 68.995 54.695 69.285 54.865 ;
        RECT 69.455 54.695 69.745 54.865 ;
        RECT 69.915 54.695 70.205 54.865 ;
        RECT 70.375 54.695 70.665 54.865 ;
        RECT 70.835 54.695 71.125 54.865 ;
        RECT 71.295 54.695 71.585 54.865 ;
        RECT 71.755 54.695 72.045 54.865 ;
        RECT 72.215 54.695 72.505 54.865 ;
        RECT 72.675 54.695 72.965 54.865 ;
        RECT 73.135 54.695 73.425 54.865 ;
        RECT 73.595 54.695 73.885 54.865 ;
        RECT 74.055 54.695 74.345 54.865 ;
        RECT 74.515 54.695 74.805 54.865 ;
        RECT 74.975 54.695 75.265 54.865 ;
        RECT 75.435 54.695 75.725 54.865 ;
        RECT 75.895 54.695 76.185 54.865 ;
        RECT 76.355 54.695 76.645 54.865 ;
        RECT 76.815 54.695 77.105 54.865 ;
        RECT 77.275 54.695 77.565 54.865 ;
        RECT 77.735 54.695 78.025 54.865 ;
        RECT 78.195 54.695 78.485 54.865 ;
        RECT 78.655 54.695 78.945 54.865 ;
        RECT 79.115 54.695 79.405 54.865 ;
        RECT 79.575 54.695 79.865 54.865 ;
        RECT 80.035 54.695 80.325 54.865 ;
        RECT 80.495 54.695 80.785 54.865 ;
        RECT 80.955 54.695 81.245 54.865 ;
        RECT 81.415 54.695 81.705 54.865 ;
        RECT 81.875 54.695 82.165 54.865 ;
        RECT 82.335 54.695 82.625 54.865 ;
        RECT 82.795 54.695 83.085 54.865 ;
        RECT 83.255 54.695 83.545 54.865 ;
        RECT 83.715 54.695 84.005 54.865 ;
        RECT 84.175 54.695 84.465 54.865 ;
        RECT 84.635 54.695 84.925 54.865 ;
        RECT 85.095 54.695 85.385 54.865 ;
        RECT 85.555 54.695 85.845 54.865 ;
        RECT 86.015 54.695 86.305 54.865 ;
        RECT 86.475 54.695 86.765 54.865 ;
        RECT 86.935 54.695 87.225 54.865 ;
        RECT 87.395 54.695 87.685 54.865 ;
        RECT 87.855 54.695 88.145 54.865 ;
        RECT 88.315 54.695 88.605 54.865 ;
        RECT 88.775 54.695 89.065 54.865 ;
        RECT 89.235 54.695 89.525 54.865 ;
        RECT 89.695 54.695 89.985 54.865 ;
        RECT 90.155 54.695 90.445 54.865 ;
        RECT 90.615 54.695 90.905 54.865 ;
        RECT 91.075 54.695 91.365 54.865 ;
        RECT 91.535 54.695 91.825 54.865 ;
        RECT 91.995 54.695 92.285 54.865 ;
        RECT 92.455 54.695 92.745 54.865 ;
        RECT 92.915 54.695 93.205 54.865 ;
        RECT 93.375 54.695 93.665 54.865 ;
        RECT 93.835 54.695 94.125 54.865 ;
        RECT 94.295 54.695 94.585 54.865 ;
        RECT 94.755 54.695 95.045 54.865 ;
        RECT 95.215 54.695 95.505 54.865 ;
        RECT 95.675 54.695 95.965 54.865 ;
        RECT 96.135 54.695 96.425 54.865 ;
        RECT 96.595 54.695 96.885 54.865 ;
        RECT 97.055 54.695 97.345 54.865 ;
        RECT 97.515 54.695 97.805 54.865 ;
        RECT 97.975 54.695 98.265 54.865 ;
        RECT 98.435 54.695 98.725 54.865 ;
        RECT 98.895 54.695 99.185 54.865 ;
        RECT 99.355 54.695 99.645 54.865 ;
        RECT 99.815 54.695 99.960 54.865 ;
        RECT 16.785 53.605 17.995 54.695 ;
        RECT 18.165 53.605 23.510 54.695 ;
        RECT 23.685 53.605 29.030 54.695 ;
        RECT 29.205 53.605 34.550 54.695 ;
        RECT 34.725 53.605 40.070 54.695 ;
        RECT 40.245 53.605 43.755 54.695 ;
        RECT 16.785 52.895 17.305 53.435 ;
        RECT 17.475 53.065 17.995 53.605 ;
        RECT 18.165 52.915 20.745 53.435 ;
        RECT 20.915 53.085 23.510 53.605 ;
        RECT 23.685 52.915 26.265 53.435 ;
        RECT 26.435 53.085 29.030 53.605 ;
        RECT 29.205 52.915 31.785 53.435 ;
        RECT 31.955 53.085 34.550 53.605 ;
        RECT 34.725 52.915 37.305 53.435 ;
        RECT 37.475 53.085 40.070 53.605 ;
        RECT 40.245 52.915 41.895 53.435 ;
        RECT 42.065 53.085 43.755 53.605 ;
        RECT 44.845 53.530 45.135 54.695 ;
        RECT 45.305 53.605 50.650 54.695 ;
        RECT 50.825 53.605 56.170 54.695 ;
        RECT 56.355 53.885 56.650 54.695 ;
        RECT 45.305 52.915 47.885 53.435 ;
        RECT 48.055 53.085 50.650 53.605 ;
        RECT 50.825 52.915 53.405 53.435 ;
        RECT 53.575 53.085 56.170 53.605 ;
        RECT 56.830 53.385 57.075 54.525 ;
        RECT 57.250 53.885 57.510 54.695 ;
        RECT 58.110 54.690 64.385 54.695 ;
        RECT 57.690 53.385 57.940 54.520 ;
        RECT 58.110 53.895 58.370 54.690 ;
      LAYER li1 ;
        RECT 58.540 53.795 58.800 54.520 ;
      LAYER li1 ;
        RECT 58.970 53.965 59.230 54.690 ;
      LAYER li1 ;
        RECT 59.400 53.795 59.660 54.520 ;
      LAYER li1 ;
        RECT 59.830 53.965 60.090 54.690 ;
      LAYER li1 ;
        RECT 60.260 53.795 60.520 54.520 ;
      LAYER li1 ;
        RECT 60.690 53.965 60.950 54.690 ;
      LAYER li1 ;
        RECT 61.120 53.795 61.380 54.520 ;
      LAYER li1 ;
        RECT 61.550 53.965 61.795 54.690 ;
      LAYER li1 ;
        RECT 61.965 53.795 62.225 54.520 ;
      LAYER li1 ;
        RECT 62.410 53.965 62.655 54.690 ;
      LAYER li1 ;
        RECT 62.825 53.795 63.085 54.520 ;
      LAYER li1 ;
        RECT 63.270 53.965 63.515 54.690 ;
      LAYER li1 ;
        RECT 63.685 53.795 63.945 54.520 ;
      LAYER li1 ;
        RECT 64.130 53.965 64.385 54.690 ;
      LAYER li1 ;
        RECT 58.540 53.780 63.945 53.795 ;
        RECT 64.555 53.780 64.845 54.520 ;
      LAYER li1 ;
        RECT 65.015 53.950 65.285 54.695 ;
      LAYER li1 ;
        RECT 58.540 53.555 65.285 53.780 ;
      LAYER li1 ;
        RECT 65.545 53.605 70.890 54.695 ;
        RECT 71.065 53.605 72.735 54.695 ;
        RECT 56.830 53.135 63.950 53.385 ;
        RECT 16.785 52.145 17.995 52.895 ;
        RECT 18.165 52.145 23.510 52.915 ;
        RECT 23.685 52.145 29.030 52.915 ;
        RECT 29.205 52.145 34.550 52.915 ;
        RECT 34.725 52.145 40.070 52.915 ;
        RECT 40.245 52.145 43.755 52.915 ;
        RECT 44.845 52.145 45.135 52.870 ;
        RECT 45.305 52.145 50.650 52.915 ;
        RECT 50.825 52.145 56.170 52.915 ;
        RECT 56.345 52.145 56.650 52.655 ;
        RECT 56.830 52.325 57.080 53.135 ;
        RECT 57.250 52.145 57.510 52.670 ;
        RECT 57.690 52.325 57.940 53.135 ;
      LAYER li1 ;
        RECT 64.120 52.965 65.285 53.555 ;
        RECT 58.540 52.795 65.285 52.965 ;
      LAYER li1 ;
        RECT 65.545 52.915 68.125 53.435 ;
        RECT 68.295 53.085 70.890 53.605 ;
        RECT 71.065 52.915 71.815 53.435 ;
        RECT 71.985 53.085 72.735 53.605 ;
        RECT 72.905 53.530 73.195 54.695 ;
        RECT 73.365 53.605 78.710 54.695 ;
        RECT 78.885 53.605 84.230 54.695 ;
        RECT 84.405 53.605 89.750 54.695 ;
        RECT 89.925 53.605 95.270 54.695 ;
        RECT 95.445 53.605 98.035 54.695 ;
        RECT 73.365 52.915 75.945 53.435 ;
        RECT 76.115 53.085 78.710 53.605 ;
        RECT 78.885 52.915 81.465 53.435 ;
        RECT 81.635 53.085 84.230 53.605 ;
        RECT 84.405 52.915 86.985 53.435 ;
        RECT 87.155 53.085 89.750 53.605 ;
        RECT 89.925 52.915 92.505 53.435 ;
        RECT 92.675 53.085 95.270 53.605 ;
        RECT 95.445 52.915 96.655 53.435 ;
        RECT 96.825 53.085 98.035 53.605 ;
        RECT 98.665 53.605 99.875 54.695 ;
        RECT 98.665 53.065 99.185 53.605 ;
        RECT 58.110 52.145 58.370 52.705 ;
      LAYER li1 ;
        RECT 58.540 52.340 58.800 52.795 ;
      LAYER li1 ;
        RECT 58.970 52.145 59.230 52.625 ;
      LAYER li1 ;
        RECT 59.400 52.340 59.660 52.795 ;
      LAYER li1 ;
        RECT 59.830 52.145 60.090 52.625 ;
      LAYER li1 ;
        RECT 60.260 52.340 60.520 52.795 ;
      LAYER li1 ;
        RECT 60.690 52.145 60.935 52.625 ;
      LAYER li1 ;
        RECT 61.105 52.340 61.380 52.795 ;
      LAYER li1 ;
        RECT 61.550 52.145 61.795 52.625 ;
      LAYER li1 ;
        RECT 61.965 52.340 62.225 52.795 ;
      LAYER li1 ;
        RECT 62.405 52.145 62.655 52.625 ;
      LAYER li1 ;
        RECT 62.825 52.340 63.085 52.795 ;
      LAYER li1 ;
        RECT 63.265 52.145 63.515 52.625 ;
      LAYER li1 ;
        RECT 63.685 52.340 63.945 52.795 ;
      LAYER li1 ;
        RECT 64.125 52.145 64.385 52.625 ;
      LAYER li1 ;
        RECT 64.555 52.340 64.815 52.795 ;
      LAYER li1 ;
        RECT 64.985 52.145 65.285 52.625 ;
        RECT 65.545 52.145 70.890 52.915 ;
        RECT 71.065 52.145 72.735 52.915 ;
        RECT 72.905 52.145 73.195 52.870 ;
        RECT 73.365 52.145 78.710 52.915 ;
        RECT 78.885 52.145 84.230 52.915 ;
        RECT 84.405 52.145 89.750 52.915 ;
        RECT 89.925 52.145 95.270 52.915 ;
        RECT 95.445 52.145 98.035 52.915 ;
        RECT 99.355 52.895 99.875 53.435 ;
        RECT 98.665 52.145 99.875 52.895 ;
        RECT 16.700 51.975 16.845 52.145 ;
        RECT 17.015 51.975 17.305 52.145 ;
        RECT 17.475 51.975 17.765 52.145 ;
        RECT 17.935 51.975 18.225 52.145 ;
        RECT 18.395 51.975 18.685 52.145 ;
        RECT 18.855 51.975 19.145 52.145 ;
        RECT 19.315 51.975 19.605 52.145 ;
        RECT 19.775 51.975 20.065 52.145 ;
        RECT 20.235 51.975 20.525 52.145 ;
        RECT 20.695 51.975 20.985 52.145 ;
        RECT 21.155 51.975 21.445 52.145 ;
        RECT 21.615 51.975 21.905 52.145 ;
        RECT 22.075 51.975 22.365 52.145 ;
        RECT 22.535 51.975 22.825 52.145 ;
        RECT 22.995 51.975 23.285 52.145 ;
        RECT 23.455 51.975 23.745 52.145 ;
        RECT 23.915 51.975 24.205 52.145 ;
        RECT 24.375 51.975 24.665 52.145 ;
        RECT 24.835 51.975 25.125 52.145 ;
        RECT 25.295 51.975 25.585 52.145 ;
        RECT 25.755 51.975 26.045 52.145 ;
        RECT 26.215 51.975 26.505 52.145 ;
        RECT 26.675 51.975 26.965 52.145 ;
        RECT 27.135 51.975 27.425 52.145 ;
        RECT 27.595 51.975 27.885 52.145 ;
        RECT 28.055 51.975 28.345 52.145 ;
        RECT 28.515 51.975 28.805 52.145 ;
        RECT 28.975 51.975 29.265 52.145 ;
        RECT 29.435 51.975 29.725 52.145 ;
        RECT 29.895 51.975 30.185 52.145 ;
        RECT 30.355 51.975 30.645 52.145 ;
        RECT 30.815 51.975 31.105 52.145 ;
        RECT 31.275 51.975 31.565 52.145 ;
        RECT 31.735 51.975 32.025 52.145 ;
        RECT 32.195 51.975 32.485 52.145 ;
        RECT 32.655 51.975 32.945 52.145 ;
        RECT 33.115 51.975 33.405 52.145 ;
        RECT 33.575 51.975 33.865 52.145 ;
        RECT 34.035 51.975 34.325 52.145 ;
        RECT 34.495 51.975 34.785 52.145 ;
        RECT 34.955 51.975 35.245 52.145 ;
        RECT 35.415 51.975 35.705 52.145 ;
        RECT 35.875 51.975 36.165 52.145 ;
        RECT 36.335 51.975 36.625 52.145 ;
        RECT 36.795 51.975 37.085 52.145 ;
        RECT 37.255 51.975 37.545 52.145 ;
        RECT 37.715 51.975 38.005 52.145 ;
        RECT 38.175 51.975 38.465 52.145 ;
        RECT 38.635 51.975 38.925 52.145 ;
        RECT 39.095 51.975 39.385 52.145 ;
        RECT 39.555 51.975 39.845 52.145 ;
        RECT 40.015 51.975 40.305 52.145 ;
        RECT 40.475 51.975 40.765 52.145 ;
        RECT 40.935 51.975 41.225 52.145 ;
        RECT 41.395 51.975 41.685 52.145 ;
        RECT 41.855 51.975 42.145 52.145 ;
        RECT 42.315 51.975 42.605 52.145 ;
        RECT 42.775 51.975 43.065 52.145 ;
        RECT 43.235 51.975 43.525 52.145 ;
        RECT 43.695 51.975 43.985 52.145 ;
        RECT 44.155 51.975 44.445 52.145 ;
        RECT 44.615 51.975 44.905 52.145 ;
        RECT 45.075 51.975 45.365 52.145 ;
        RECT 45.535 51.975 45.825 52.145 ;
        RECT 45.995 51.975 46.285 52.145 ;
        RECT 46.455 51.975 46.745 52.145 ;
        RECT 46.915 51.975 47.205 52.145 ;
        RECT 47.375 51.975 47.665 52.145 ;
        RECT 47.835 51.975 48.125 52.145 ;
        RECT 48.295 51.975 48.585 52.145 ;
        RECT 48.755 51.975 49.045 52.145 ;
        RECT 49.215 51.975 49.505 52.145 ;
        RECT 49.675 51.975 49.965 52.145 ;
        RECT 50.135 51.975 50.425 52.145 ;
        RECT 50.595 51.975 50.885 52.145 ;
        RECT 51.055 51.975 51.345 52.145 ;
        RECT 51.515 51.975 51.805 52.145 ;
        RECT 51.975 51.975 52.265 52.145 ;
        RECT 52.435 51.975 52.725 52.145 ;
        RECT 52.895 51.975 53.185 52.145 ;
        RECT 53.355 51.975 53.645 52.145 ;
        RECT 53.815 51.975 54.105 52.145 ;
        RECT 54.275 51.975 54.565 52.145 ;
        RECT 54.735 51.975 55.025 52.145 ;
        RECT 55.195 51.975 55.485 52.145 ;
        RECT 55.655 51.975 55.945 52.145 ;
        RECT 56.115 51.975 56.405 52.145 ;
        RECT 56.575 51.975 56.865 52.145 ;
        RECT 57.035 51.975 57.325 52.145 ;
        RECT 57.495 51.975 57.785 52.145 ;
        RECT 57.955 51.975 58.245 52.145 ;
        RECT 58.415 51.975 58.705 52.145 ;
        RECT 58.875 51.975 59.165 52.145 ;
        RECT 59.335 51.975 59.625 52.145 ;
        RECT 59.795 51.975 60.085 52.145 ;
        RECT 60.255 51.975 60.545 52.145 ;
        RECT 60.715 51.975 61.005 52.145 ;
        RECT 61.175 51.975 61.465 52.145 ;
        RECT 61.635 51.975 61.925 52.145 ;
        RECT 62.095 51.975 62.385 52.145 ;
        RECT 62.555 51.975 62.845 52.145 ;
        RECT 63.015 51.975 63.305 52.145 ;
        RECT 63.475 51.975 63.765 52.145 ;
        RECT 63.935 51.975 64.225 52.145 ;
        RECT 64.395 51.975 64.685 52.145 ;
        RECT 64.855 51.975 65.145 52.145 ;
        RECT 65.315 51.975 65.605 52.145 ;
        RECT 65.775 51.975 66.065 52.145 ;
        RECT 66.235 51.975 66.525 52.145 ;
        RECT 66.695 51.975 66.985 52.145 ;
        RECT 67.155 51.975 67.445 52.145 ;
        RECT 67.615 51.975 67.905 52.145 ;
        RECT 68.075 51.975 68.365 52.145 ;
        RECT 68.535 51.975 68.825 52.145 ;
        RECT 68.995 51.975 69.285 52.145 ;
        RECT 69.455 51.975 69.745 52.145 ;
        RECT 69.915 51.975 70.205 52.145 ;
        RECT 70.375 51.975 70.665 52.145 ;
        RECT 70.835 51.975 71.125 52.145 ;
        RECT 71.295 51.975 71.585 52.145 ;
        RECT 71.755 51.975 72.045 52.145 ;
        RECT 72.215 51.975 72.505 52.145 ;
        RECT 72.675 51.975 72.965 52.145 ;
        RECT 73.135 51.975 73.425 52.145 ;
        RECT 73.595 51.975 73.885 52.145 ;
        RECT 74.055 51.975 74.345 52.145 ;
        RECT 74.515 51.975 74.805 52.145 ;
        RECT 74.975 51.975 75.265 52.145 ;
        RECT 75.435 51.975 75.725 52.145 ;
        RECT 75.895 51.975 76.185 52.145 ;
        RECT 76.355 51.975 76.645 52.145 ;
        RECT 76.815 51.975 77.105 52.145 ;
        RECT 77.275 51.975 77.565 52.145 ;
        RECT 77.735 51.975 78.025 52.145 ;
        RECT 78.195 51.975 78.485 52.145 ;
        RECT 78.655 51.975 78.945 52.145 ;
        RECT 79.115 51.975 79.405 52.145 ;
        RECT 79.575 51.975 79.865 52.145 ;
        RECT 80.035 51.975 80.325 52.145 ;
        RECT 80.495 51.975 80.785 52.145 ;
        RECT 80.955 51.975 81.245 52.145 ;
        RECT 81.415 51.975 81.705 52.145 ;
        RECT 81.875 51.975 82.165 52.145 ;
        RECT 82.335 51.975 82.625 52.145 ;
        RECT 82.795 51.975 83.085 52.145 ;
        RECT 83.255 51.975 83.545 52.145 ;
        RECT 83.715 51.975 84.005 52.145 ;
        RECT 84.175 51.975 84.465 52.145 ;
        RECT 84.635 51.975 84.925 52.145 ;
        RECT 85.095 51.975 85.385 52.145 ;
        RECT 85.555 51.975 85.845 52.145 ;
        RECT 86.015 51.975 86.305 52.145 ;
        RECT 86.475 51.975 86.765 52.145 ;
        RECT 86.935 51.975 87.225 52.145 ;
        RECT 87.395 51.975 87.685 52.145 ;
        RECT 87.855 51.975 88.145 52.145 ;
        RECT 88.315 51.975 88.605 52.145 ;
        RECT 88.775 51.975 89.065 52.145 ;
        RECT 89.235 51.975 89.525 52.145 ;
        RECT 89.695 51.975 89.985 52.145 ;
        RECT 90.155 51.975 90.445 52.145 ;
        RECT 90.615 51.975 90.905 52.145 ;
        RECT 91.075 51.975 91.365 52.145 ;
        RECT 91.535 51.975 91.825 52.145 ;
        RECT 91.995 51.975 92.285 52.145 ;
        RECT 92.455 51.975 92.745 52.145 ;
        RECT 92.915 51.975 93.205 52.145 ;
        RECT 93.375 51.975 93.665 52.145 ;
        RECT 93.835 51.975 94.125 52.145 ;
        RECT 94.295 51.975 94.585 52.145 ;
        RECT 94.755 51.975 95.045 52.145 ;
        RECT 95.215 51.975 95.505 52.145 ;
        RECT 95.675 51.975 95.965 52.145 ;
        RECT 96.135 51.975 96.425 52.145 ;
        RECT 96.595 51.975 96.885 52.145 ;
        RECT 97.055 51.975 97.345 52.145 ;
        RECT 97.515 51.975 97.805 52.145 ;
        RECT 97.975 51.975 98.265 52.145 ;
        RECT 98.435 51.975 98.725 52.145 ;
        RECT 98.895 51.975 99.185 52.145 ;
        RECT 99.355 51.975 99.645 52.145 ;
        RECT 99.815 51.975 99.960 52.145 ;
        RECT 16.785 51.225 17.995 51.975 ;
        RECT 16.785 50.685 17.305 51.225 ;
        RECT 18.165 51.205 23.510 51.975 ;
        RECT 23.685 51.205 29.030 51.975 ;
        RECT 29.205 51.205 30.875 51.975 ;
        RECT 31.045 51.250 31.335 51.975 ;
        RECT 31.505 51.205 36.850 51.975 ;
        RECT 37.025 51.205 42.370 51.975 ;
        RECT 42.545 51.205 47.890 51.975 ;
        RECT 48.065 51.205 53.410 51.975 ;
        RECT 53.585 51.205 58.930 51.975 ;
        RECT 59.105 51.250 59.395 51.975 ;
        RECT 59.565 51.225 60.775 51.975 ;
        RECT 61.035 51.425 61.205 51.715 ;
        RECT 61.375 51.595 61.705 51.975 ;
        RECT 61.035 51.255 61.700 51.425 ;
        RECT 17.475 50.515 17.995 51.055 ;
        RECT 18.165 50.685 20.745 51.205 ;
        RECT 20.915 50.515 23.510 51.035 ;
        RECT 23.685 50.685 26.265 51.205 ;
        RECT 26.435 50.515 29.030 51.035 ;
        RECT 29.205 50.685 29.955 51.205 ;
        RECT 30.125 50.515 30.875 51.035 ;
        RECT 31.505 50.685 34.085 51.205 ;
        RECT 16.785 49.425 17.995 50.515 ;
        RECT 18.165 49.425 23.510 50.515 ;
        RECT 23.685 49.425 29.030 50.515 ;
        RECT 29.205 49.425 30.875 50.515 ;
        RECT 31.045 49.425 31.335 50.590 ;
        RECT 34.255 50.515 36.850 51.035 ;
        RECT 37.025 50.685 39.605 51.205 ;
        RECT 39.775 50.515 42.370 51.035 ;
        RECT 42.545 50.685 45.125 51.205 ;
        RECT 45.295 50.515 47.890 51.035 ;
        RECT 48.065 50.685 50.645 51.205 ;
        RECT 50.815 50.515 53.410 51.035 ;
        RECT 53.585 50.685 56.165 51.205 ;
        RECT 56.335 50.515 58.930 51.035 ;
        RECT 59.565 50.685 60.085 51.225 ;
        RECT 31.505 49.425 36.850 50.515 ;
        RECT 37.025 49.425 42.370 50.515 ;
        RECT 42.545 49.425 47.890 50.515 ;
        RECT 48.065 49.425 53.410 50.515 ;
        RECT 53.585 49.425 58.930 50.515 ;
        RECT 59.105 49.425 59.395 50.590 ;
        RECT 60.255 50.515 60.775 51.055 ;
        RECT 59.565 49.425 60.775 50.515 ;
      LAYER li1 ;
        RECT 60.950 50.435 61.300 51.085 ;
      LAYER li1 ;
        RECT 61.470 50.265 61.700 51.255 ;
        RECT 61.035 50.095 61.700 50.265 ;
        RECT 61.035 49.595 61.205 50.095 ;
        RECT 61.375 49.425 61.705 49.925 ;
        RECT 61.875 49.595 62.100 51.715 ;
        RECT 62.315 51.515 62.565 51.975 ;
        RECT 62.750 51.525 63.080 51.695 ;
        RECT 63.260 51.525 64.010 51.695 ;
      LAYER li1 ;
        RECT 62.300 50.395 62.580 50.995 ;
      LAYER li1 ;
        RECT 62.750 49.995 62.920 51.525 ;
        RECT 63.090 51.025 63.670 51.355 ;
        RECT 63.090 50.155 63.330 51.025 ;
        RECT 63.840 50.745 64.010 51.525 ;
        RECT 64.260 51.475 64.630 51.975 ;
        RECT 64.810 51.525 65.270 51.695 ;
        RECT 65.500 51.525 66.170 51.695 ;
        RECT 64.810 51.295 64.980 51.525 ;
        RECT 64.180 50.995 64.980 51.295 ;
        RECT 65.150 51.025 65.700 51.355 ;
        RECT 64.180 50.965 64.350 50.995 ;
        RECT 64.470 50.745 64.640 50.815 ;
        RECT 63.840 50.575 64.640 50.745 ;
        RECT 64.130 50.485 64.640 50.575 ;
        RECT 63.520 50.050 63.960 50.405 ;
        RECT 62.300 49.425 62.565 49.885 ;
        RECT 62.750 49.620 62.985 49.995 ;
        RECT 64.130 49.870 64.300 50.485 ;
        RECT 63.230 49.700 64.300 49.870 ;
        RECT 64.470 49.425 64.640 50.225 ;
        RECT 64.810 49.925 64.980 50.995 ;
        RECT 65.150 50.095 65.340 50.815 ;
        RECT 65.510 50.485 65.700 51.025 ;
        RECT 66.000 50.985 66.170 51.525 ;
        RECT 66.485 51.445 66.655 51.975 ;
        RECT 66.950 51.325 67.310 51.765 ;
        RECT 67.485 51.495 67.655 51.975 ;
        RECT 68.355 51.500 68.525 51.975 ;
        RECT 69.205 51.500 69.375 51.975 ;
        RECT 66.950 51.155 67.450 51.325 ;
        RECT 67.280 50.985 67.450 51.155 ;
        RECT 69.685 51.205 75.030 51.975 ;
        RECT 75.205 51.205 80.550 51.975 ;
        RECT 80.725 51.205 86.070 51.975 ;
        RECT 87.165 51.250 87.455 51.975 ;
        RECT 87.625 51.205 92.970 51.975 ;
        RECT 93.145 51.205 98.490 51.975 ;
        RECT 98.665 51.225 99.875 51.975 ;
        RECT 66.000 50.815 67.090 50.985 ;
        RECT 67.280 50.815 69.100 50.985 ;
        RECT 65.510 50.155 65.830 50.485 ;
        RECT 64.810 49.595 65.060 49.925 ;
        RECT 66.000 49.895 66.170 50.815 ;
        RECT 67.280 50.560 67.450 50.815 ;
        RECT 69.685 50.685 72.265 51.205 ;
        RECT 66.340 50.390 67.450 50.560 ;
        RECT 72.435 50.515 75.030 51.035 ;
        RECT 75.205 50.685 77.785 51.205 ;
        RECT 77.955 50.515 80.550 51.035 ;
        RECT 80.725 50.685 83.305 51.205 ;
        RECT 83.475 50.515 86.070 51.035 ;
        RECT 87.625 50.685 90.205 51.205 ;
        RECT 66.340 50.230 67.200 50.390 ;
        RECT 65.285 49.725 66.170 49.895 ;
        RECT 66.350 49.425 66.565 49.925 ;
        RECT 67.030 49.605 67.200 50.230 ;
        RECT 67.485 49.425 67.665 50.205 ;
        RECT 68.360 49.425 68.530 50.255 ;
        RECT 69.200 49.425 69.370 50.255 ;
        RECT 69.685 49.425 75.030 50.515 ;
        RECT 75.205 49.425 80.550 50.515 ;
        RECT 80.725 49.425 86.070 50.515 ;
        RECT 87.165 49.425 87.455 50.590 ;
        RECT 90.375 50.515 92.970 51.035 ;
        RECT 93.145 50.685 95.725 51.205 ;
        RECT 95.895 50.515 98.490 51.035 ;
        RECT 87.625 49.425 92.970 50.515 ;
        RECT 93.145 49.425 98.490 50.515 ;
        RECT 98.665 50.515 99.185 51.055 ;
        RECT 99.355 50.685 99.875 51.225 ;
        RECT 98.665 49.425 99.875 50.515 ;
        RECT 16.700 49.255 16.845 49.425 ;
        RECT 17.015 49.255 17.305 49.425 ;
        RECT 17.475 49.255 17.765 49.425 ;
        RECT 17.935 49.255 18.225 49.425 ;
        RECT 18.395 49.255 18.685 49.425 ;
        RECT 18.855 49.255 19.145 49.425 ;
        RECT 19.315 49.255 19.605 49.425 ;
        RECT 19.775 49.255 20.065 49.425 ;
        RECT 20.235 49.255 20.525 49.425 ;
        RECT 20.695 49.255 20.985 49.425 ;
        RECT 21.155 49.255 21.445 49.425 ;
        RECT 21.615 49.255 21.905 49.425 ;
        RECT 22.075 49.255 22.365 49.425 ;
        RECT 22.535 49.255 22.825 49.425 ;
        RECT 22.995 49.255 23.285 49.425 ;
        RECT 23.455 49.255 23.745 49.425 ;
        RECT 23.915 49.255 24.205 49.425 ;
        RECT 24.375 49.255 24.665 49.425 ;
        RECT 24.835 49.255 25.125 49.425 ;
        RECT 25.295 49.255 25.585 49.425 ;
        RECT 25.755 49.255 26.045 49.425 ;
        RECT 26.215 49.255 26.505 49.425 ;
        RECT 26.675 49.255 26.965 49.425 ;
        RECT 27.135 49.255 27.425 49.425 ;
        RECT 27.595 49.255 27.885 49.425 ;
        RECT 28.055 49.255 28.345 49.425 ;
        RECT 28.515 49.255 28.805 49.425 ;
        RECT 28.975 49.255 29.265 49.425 ;
        RECT 29.435 49.255 29.725 49.425 ;
        RECT 29.895 49.255 30.185 49.425 ;
        RECT 30.355 49.255 30.645 49.425 ;
        RECT 30.815 49.255 31.105 49.425 ;
        RECT 31.275 49.255 31.565 49.425 ;
        RECT 31.735 49.255 32.025 49.425 ;
        RECT 32.195 49.255 32.485 49.425 ;
        RECT 32.655 49.255 32.945 49.425 ;
        RECT 33.115 49.255 33.405 49.425 ;
        RECT 33.575 49.255 33.865 49.425 ;
        RECT 34.035 49.255 34.325 49.425 ;
        RECT 34.495 49.255 34.785 49.425 ;
        RECT 34.955 49.255 35.245 49.425 ;
        RECT 35.415 49.255 35.705 49.425 ;
        RECT 35.875 49.255 36.165 49.425 ;
        RECT 36.335 49.255 36.625 49.425 ;
        RECT 36.795 49.255 37.085 49.425 ;
        RECT 37.255 49.255 37.545 49.425 ;
        RECT 37.715 49.255 38.005 49.425 ;
        RECT 38.175 49.255 38.465 49.425 ;
        RECT 38.635 49.255 38.925 49.425 ;
        RECT 39.095 49.255 39.385 49.425 ;
        RECT 39.555 49.255 39.845 49.425 ;
        RECT 40.015 49.255 40.305 49.425 ;
        RECT 40.475 49.255 40.765 49.425 ;
        RECT 40.935 49.255 41.225 49.425 ;
        RECT 41.395 49.255 41.685 49.425 ;
        RECT 41.855 49.255 42.145 49.425 ;
        RECT 42.315 49.255 42.605 49.425 ;
        RECT 42.775 49.255 43.065 49.425 ;
        RECT 43.235 49.255 43.525 49.425 ;
        RECT 43.695 49.255 43.985 49.425 ;
        RECT 44.155 49.255 44.445 49.425 ;
        RECT 44.615 49.255 44.905 49.425 ;
        RECT 45.075 49.255 45.365 49.425 ;
        RECT 45.535 49.255 45.825 49.425 ;
        RECT 45.995 49.255 46.285 49.425 ;
        RECT 46.455 49.255 46.745 49.425 ;
        RECT 46.915 49.255 47.205 49.425 ;
        RECT 47.375 49.255 47.665 49.425 ;
        RECT 47.835 49.255 48.125 49.425 ;
        RECT 48.295 49.255 48.585 49.425 ;
        RECT 48.755 49.255 49.045 49.425 ;
        RECT 49.215 49.255 49.505 49.425 ;
        RECT 49.675 49.255 49.965 49.425 ;
        RECT 50.135 49.255 50.425 49.425 ;
        RECT 50.595 49.255 50.885 49.425 ;
        RECT 51.055 49.255 51.345 49.425 ;
        RECT 51.515 49.255 51.805 49.425 ;
        RECT 51.975 49.255 52.265 49.425 ;
        RECT 52.435 49.255 52.725 49.425 ;
        RECT 52.895 49.255 53.185 49.425 ;
        RECT 53.355 49.255 53.645 49.425 ;
        RECT 53.815 49.255 54.105 49.425 ;
        RECT 54.275 49.255 54.565 49.425 ;
        RECT 54.735 49.255 55.025 49.425 ;
        RECT 55.195 49.255 55.485 49.425 ;
        RECT 55.655 49.255 55.945 49.425 ;
        RECT 56.115 49.255 56.405 49.425 ;
        RECT 56.575 49.255 56.865 49.425 ;
        RECT 57.035 49.255 57.325 49.425 ;
        RECT 57.495 49.255 57.785 49.425 ;
        RECT 57.955 49.255 58.245 49.425 ;
        RECT 58.415 49.255 58.705 49.425 ;
        RECT 58.875 49.255 59.165 49.425 ;
        RECT 59.335 49.255 59.625 49.425 ;
        RECT 59.795 49.255 60.085 49.425 ;
        RECT 60.255 49.255 60.545 49.425 ;
        RECT 60.715 49.255 61.005 49.425 ;
        RECT 61.175 49.255 61.465 49.425 ;
        RECT 61.635 49.255 61.925 49.425 ;
        RECT 62.095 49.255 62.385 49.425 ;
        RECT 62.555 49.255 62.845 49.425 ;
        RECT 63.015 49.255 63.305 49.425 ;
        RECT 63.475 49.255 63.765 49.425 ;
        RECT 63.935 49.255 64.225 49.425 ;
        RECT 64.395 49.255 64.685 49.425 ;
        RECT 64.855 49.255 65.145 49.425 ;
        RECT 65.315 49.255 65.605 49.425 ;
        RECT 65.775 49.255 66.065 49.425 ;
        RECT 66.235 49.255 66.525 49.425 ;
        RECT 66.695 49.255 66.985 49.425 ;
        RECT 67.155 49.255 67.445 49.425 ;
        RECT 67.615 49.255 67.905 49.425 ;
        RECT 68.075 49.255 68.365 49.425 ;
        RECT 68.535 49.255 68.825 49.425 ;
        RECT 68.995 49.255 69.285 49.425 ;
        RECT 69.455 49.255 69.745 49.425 ;
        RECT 69.915 49.255 70.205 49.425 ;
        RECT 70.375 49.255 70.665 49.425 ;
        RECT 70.835 49.255 71.125 49.425 ;
        RECT 71.295 49.255 71.585 49.425 ;
        RECT 71.755 49.255 72.045 49.425 ;
        RECT 72.215 49.255 72.505 49.425 ;
        RECT 72.675 49.255 72.965 49.425 ;
        RECT 73.135 49.255 73.425 49.425 ;
        RECT 73.595 49.255 73.885 49.425 ;
        RECT 74.055 49.255 74.345 49.425 ;
        RECT 74.515 49.255 74.805 49.425 ;
        RECT 74.975 49.255 75.265 49.425 ;
        RECT 75.435 49.255 75.725 49.425 ;
        RECT 75.895 49.255 76.185 49.425 ;
        RECT 76.355 49.255 76.645 49.425 ;
        RECT 76.815 49.255 77.105 49.425 ;
        RECT 77.275 49.255 77.565 49.425 ;
        RECT 77.735 49.255 78.025 49.425 ;
        RECT 78.195 49.255 78.485 49.425 ;
        RECT 78.655 49.255 78.945 49.425 ;
        RECT 79.115 49.255 79.405 49.425 ;
        RECT 79.575 49.255 79.865 49.425 ;
        RECT 80.035 49.255 80.325 49.425 ;
        RECT 80.495 49.255 80.785 49.425 ;
        RECT 80.955 49.255 81.245 49.425 ;
        RECT 81.415 49.255 81.705 49.425 ;
        RECT 81.875 49.255 82.165 49.425 ;
        RECT 82.335 49.255 82.625 49.425 ;
        RECT 82.795 49.255 83.085 49.425 ;
        RECT 83.255 49.255 83.545 49.425 ;
        RECT 83.715 49.255 84.005 49.425 ;
        RECT 84.175 49.255 84.465 49.425 ;
        RECT 84.635 49.255 84.925 49.425 ;
        RECT 85.095 49.255 85.385 49.425 ;
        RECT 85.555 49.255 85.845 49.425 ;
        RECT 86.015 49.255 86.305 49.425 ;
        RECT 86.475 49.255 86.765 49.425 ;
        RECT 86.935 49.255 87.225 49.425 ;
        RECT 87.395 49.255 87.685 49.425 ;
        RECT 87.855 49.255 88.145 49.425 ;
        RECT 88.315 49.255 88.605 49.425 ;
        RECT 88.775 49.255 89.065 49.425 ;
        RECT 89.235 49.255 89.525 49.425 ;
        RECT 89.695 49.255 89.985 49.425 ;
        RECT 90.155 49.255 90.445 49.425 ;
        RECT 90.615 49.255 90.905 49.425 ;
        RECT 91.075 49.255 91.365 49.425 ;
        RECT 91.535 49.255 91.825 49.425 ;
        RECT 91.995 49.255 92.285 49.425 ;
        RECT 92.455 49.255 92.745 49.425 ;
        RECT 92.915 49.255 93.205 49.425 ;
        RECT 93.375 49.255 93.665 49.425 ;
        RECT 93.835 49.255 94.125 49.425 ;
        RECT 94.295 49.255 94.585 49.425 ;
        RECT 94.755 49.255 95.045 49.425 ;
        RECT 95.215 49.255 95.505 49.425 ;
        RECT 95.675 49.255 95.965 49.425 ;
        RECT 96.135 49.255 96.425 49.425 ;
        RECT 96.595 49.255 96.885 49.425 ;
        RECT 97.055 49.255 97.345 49.425 ;
        RECT 97.515 49.255 97.805 49.425 ;
        RECT 97.975 49.255 98.265 49.425 ;
        RECT 98.435 49.255 98.725 49.425 ;
        RECT 98.895 49.255 99.185 49.425 ;
        RECT 99.355 49.255 99.645 49.425 ;
        RECT 99.815 49.255 99.960 49.425 ;
        RECT 16.785 48.165 17.995 49.255 ;
        RECT 18.165 48.165 19.375 49.255 ;
        RECT 19.735 48.530 20.065 49.255 ;
        RECT 16.785 47.455 17.305 47.995 ;
        RECT 17.475 47.625 17.995 48.165 ;
        RECT 18.165 47.455 18.685 47.995 ;
        RECT 18.855 47.625 19.375 48.165 ;
        RECT 16.785 46.705 17.995 47.455 ;
        RECT 18.165 46.705 19.375 47.455 ;
      LAYER li1 ;
        RECT 19.545 46.875 20.065 48.360 ;
      LAYER li1 ;
        RECT 20.925 48.165 26.270 49.255 ;
        RECT 26.445 48.165 31.790 49.255 ;
        RECT 31.965 48.165 37.310 49.255 ;
        RECT 37.485 48.165 42.830 49.255 ;
        RECT 43.005 48.165 44.675 49.255 ;
        RECT 20.925 47.475 23.505 47.995 ;
        RECT 23.675 47.645 26.270 48.165 ;
        RECT 26.445 47.475 29.025 47.995 ;
        RECT 29.195 47.645 31.790 48.165 ;
        RECT 31.965 47.475 34.545 47.995 ;
        RECT 34.715 47.645 37.310 48.165 ;
        RECT 37.485 47.475 40.065 47.995 ;
        RECT 40.235 47.645 42.830 48.165 ;
        RECT 43.005 47.475 43.755 47.995 ;
        RECT 43.925 47.645 44.675 48.165 ;
        RECT 44.845 48.090 45.135 49.255 ;
        RECT 45.305 48.165 50.650 49.255 ;
        RECT 50.825 48.165 56.170 49.255 ;
        RECT 56.345 48.165 58.935 49.255 ;
        RECT 45.305 47.475 47.885 47.995 ;
        RECT 48.055 47.645 50.650 48.165 ;
        RECT 50.825 47.475 53.405 47.995 ;
        RECT 53.575 47.645 56.170 48.165 ;
        RECT 56.345 47.475 57.555 47.995 ;
        RECT 57.725 47.645 58.935 48.165 ;
      LAYER li1 ;
        RECT 59.565 48.180 59.835 49.085 ;
      LAYER li1 ;
        RECT 60.005 48.495 60.335 49.255 ;
        RECT 60.515 48.325 60.685 49.085 ;
        RECT 20.235 46.705 20.575 47.365 ;
        RECT 20.925 46.705 26.270 47.475 ;
        RECT 26.445 46.705 31.790 47.475 ;
        RECT 31.965 46.705 37.310 47.475 ;
        RECT 37.485 46.705 42.830 47.475 ;
        RECT 43.005 46.705 44.675 47.475 ;
        RECT 44.845 46.705 45.135 47.430 ;
        RECT 45.305 46.705 50.650 47.475 ;
        RECT 50.825 46.705 56.170 47.475 ;
        RECT 56.345 46.705 58.935 47.475 ;
      LAYER li1 ;
        RECT 59.565 47.380 59.735 48.180 ;
      LAYER li1 ;
        RECT 60.020 48.155 60.685 48.325 ;
        RECT 60.945 48.165 66.290 49.255 ;
        RECT 66.465 48.165 71.810 49.255 ;
        RECT 60.020 48.010 60.190 48.155 ;
        RECT 59.905 47.680 60.190 48.010 ;
        RECT 60.020 47.425 60.190 47.680 ;
      LAYER li1 ;
        RECT 60.425 47.605 60.755 47.975 ;
      LAYER li1 ;
        RECT 60.945 47.475 63.525 47.995 ;
        RECT 63.695 47.645 66.290 48.165 ;
        RECT 66.465 47.475 69.045 47.995 ;
        RECT 69.215 47.645 71.810 48.165 ;
        RECT 72.905 48.090 73.195 49.255 ;
        RECT 73.365 48.165 78.710 49.255 ;
        RECT 78.885 48.165 84.230 49.255 ;
        RECT 84.405 48.165 89.750 49.255 ;
        RECT 89.925 48.165 95.270 49.255 ;
        RECT 95.445 48.165 98.035 49.255 ;
        RECT 73.365 47.475 75.945 47.995 ;
        RECT 76.115 47.645 78.710 48.165 ;
        RECT 78.885 47.475 81.465 47.995 ;
        RECT 81.635 47.645 84.230 48.165 ;
        RECT 84.405 47.475 86.985 47.995 ;
        RECT 87.155 47.645 89.750 48.165 ;
        RECT 89.925 47.475 92.505 47.995 ;
        RECT 92.675 47.645 95.270 48.165 ;
        RECT 95.445 47.475 96.655 47.995 ;
        RECT 96.825 47.645 98.035 48.165 ;
        RECT 98.665 48.165 99.875 49.255 ;
        RECT 98.665 47.625 99.185 48.165 ;
      LAYER li1 ;
        RECT 59.565 46.875 59.825 47.380 ;
      LAYER li1 ;
        RECT 60.020 47.255 60.685 47.425 ;
        RECT 60.005 46.705 60.335 47.085 ;
        RECT 60.515 46.875 60.685 47.255 ;
        RECT 60.945 46.705 66.290 47.475 ;
        RECT 66.465 46.705 71.810 47.475 ;
        RECT 72.905 46.705 73.195 47.430 ;
        RECT 73.365 46.705 78.710 47.475 ;
        RECT 78.885 46.705 84.230 47.475 ;
        RECT 84.405 46.705 89.750 47.475 ;
        RECT 89.925 46.705 95.270 47.475 ;
        RECT 95.445 46.705 98.035 47.475 ;
        RECT 99.355 47.455 99.875 47.995 ;
        RECT 98.665 46.705 99.875 47.455 ;
        RECT 16.700 46.535 16.845 46.705 ;
        RECT 17.015 46.535 17.305 46.705 ;
        RECT 17.475 46.535 17.765 46.705 ;
        RECT 17.935 46.535 18.225 46.705 ;
        RECT 18.395 46.535 18.685 46.705 ;
        RECT 18.855 46.535 19.145 46.705 ;
        RECT 19.315 46.535 19.605 46.705 ;
        RECT 19.775 46.535 20.065 46.705 ;
        RECT 20.235 46.535 20.525 46.705 ;
        RECT 20.695 46.535 20.985 46.705 ;
        RECT 21.155 46.535 21.445 46.705 ;
        RECT 21.615 46.535 21.905 46.705 ;
        RECT 22.075 46.535 22.365 46.705 ;
        RECT 22.535 46.535 22.825 46.705 ;
        RECT 22.995 46.535 23.285 46.705 ;
        RECT 23.455 46.535 23.745 46.705 ;
        RECT 23.915 46.535 24.205 46.705 ;
        RECT 24.375 46.535 24.665 46.705 ;
        RECT 24.835 46.535 25.125 46.705 ;
        RECT 25.295 46.535 25.585 46.705 ;
        RECT 25.755 46.535 26.045 46.705 ;
        RECT 26.215 46.535 26.505 46.705 ;
        RECT 26.675 46.535 26.965 46.705 ;
        RECT 27.135 46.535 27.425 46.705 ;
        RECT 27.595 46.535 27.885 46.705 ;
        RECT 28.055 46.535 28.345 46.705 ;
        RECT 28.515 46.535 28.805 46.705 ;
        RECT 28.975 46.535 29.265 46.705 ;
        RECT 29.435 46.535 29.725 46.705 ;
        RECT 29.895 46.535 30.185 46.705 ;
        RECT 30.355 46.535 30.645 46.705 ;
        RECT 30.815 46.535 31.105 46.705 ;
        RECT 31.275 46.535 31.565 46.705 ;
        RECT 31.735 46.535 32.025 46.705 ;
        RECT 32.195 46.535 32.485 46.705 ;
        RECT 32.655 46.535 32.945 46.705 ;
        RECT 33.115 46.535 33.405 46.705 ;
        RECT 33.575 46.535 33.865 46.705 ;
        RECT 34.035 46.535 34.325 46.705 ;
        RECT 34.495 46.535 34.785 46.705 ;
        RECT 34.955 46.535 35.245 46.705 ;
        RECT 35.415 46.535 35.705 46.705 ;
        RECT 35.875 46.535 36.165 46.705 ;
        RECT 36.335 46.535 36.625 46.705 ;
        RECT 36.795 46.535 37.085 46.705 ;
        RECT 37.255 46.535 37.545 46.705 ;
        RECT 37.715 46.535 38.005 46.705 ;
        RECT 38.175 46.535 38.465 46.705 ;
        RECT 38.635 46.535 38.925 46.705 ;
        RECT 39.095 46.535 39.385 46.705 ;
        RECT 39.555 46.535 39.845 46.705 ;
        RECT 40.015 46.535 40.305 46.705 ;
        RECT 40.475 46.535 40.765 46.705 ;
        RECT 40.935 46.535 41.225 46.705 ;
        RECT 41.395 46.535 41.685 46.705 ;
        RECT 41.855 46.535 42.145 46.705 ;
        RECT 42.315 46.535 42.605 46.705 ;
        RECT 42.775 46.535 43.065 46.705 ;
        RECT 43.235 46.535 43.525 46.705 ;
        RECT 43.695 46.535 43.985 46.705 ;
        RECT 44.155 46.535 44.445 46.705 ;
        RECT 44.615 46.535 44.905 46.705 ;
        RECT 45.075 46.535 45.365 46.705 ;
        RECT 45.535 46.535 45.825 46.705 ;
        RECT 45.995 46.535 46.285 46.705 ;
        RECT 46.455 46.535 46.745 46.705 ;
        RECT 46.915 46.535 47.205 46.705 ;
        RECT 47.375 46.535 47.665 46.705 ;
        RECT 47.835 46.535 48.125 46.705 ;
        RECT 48.295 46.535 48.585 46.705 ;
        RECT 48.755 46.535 49.045 46.705 ;
        RECT 49.215 46.535 49.505 46.705 ;
        RECT 49.675 46.535 49.965 46.705 ;
        RECT 50.135 46.535 50.425 46.705 ;
        RECT 50.595 46.535 50.885 46.705 ;
        RECT 51.055 46.535 51.345 46.705 ;
        RECT 51.515 46.535 51.805 46.705 ;
        RECT 51.975 46.535 52.265 46.705 ;
        RECT 52.435 46.535 52.725 46.705 ;
        RECT 52.895 46.535 53.185 46.705 ;
        RECT 53.355 46.535 53.645 46.705 ;
        RECT 53.815 46.535 54.105 46.705 ;
        RECT 54.275 46.535 54.565 46.705 ;
        RECT 54.735 46.535 55.025 46.705 ;
        RECT 55.195 46.535 55.485 46.705 ;
        RECT 55.655 46.535 55.945 46.705 ;
        RECT 56.115 46.535 56.405 46.705 ;
        RECT 56.575 46.535 56.865 46.705 ;
        RECT 57.035 46.535 57.325 46.705 ;
        RECT 57.495 46.535 57.785 46.705 ;
        RECT 57.955 46.535 58.245 46.705 ;
        RECT 58.415 46.535 58.705 46.705 ;
        RECT 58.875 46.535 59.165 46.705 ;
        RECT 59.335 46.535 59.625 46.705 ;
        RECT 59.795 46.535 60.085 46.705 ;
        RECT 60.255 46.535 60.545 46.705 ;
        RECT 60.715 46.535 61.005 46.705 ;
        RECT 61.175 46.535 61.465 46.705 ;
        RECT 61.635 46.535 61.925 46.705 ;
        RECT 62.095 46.535 62.385 46.705 ;
        RECT 62.555 46.535 62.845 46.705 ;
        RECT 63.015 46.535 63.305 46.705 ;
        RECT 63.475 46.535 63.765 46.705 ;
        RECT 63.935 46.535 64.225 46.705 ;
        RECT 64.395 46.535 64.685 46.705 ;
        RECT 64.855 46.535 65.145 46.705 ;
        RECT 65.315 46.535 65.605 46.705 ;
        RECT 65.775 46.535 66.065 46.705 ;
        RECT 66.235 46.535 66.525 46.705 ;
        RECT 66.695 46.535 66.985 46.705 ;
        RECT 67.155 46.535 67.445 46.705 ;
        RECT 67.615 46.535 67.905 46.705 ;
        RECT 68.075 46.535 68.365 46.705 ;
        RECT 68.535 46.535 68.825 46.705 ;
        RECT 68.995 46.535 69.285 46.705 ;
        RECT 69.455 46.535 69.745 46.705 ;
        RECT 69.915 46.535 70.205 46.705 ;
        RECT 70.375 46.535 70.665 46.705 ;
        RECT 70.835 46.535 71.125 46.705 ;
        RECT 71.295 46.535 71.585 46.705 ;
        RECT 71.755 46.535 72.045 46.705 ;
        RECT 72.215 46.535 72.505 46.705 ;
        RECT 72.675 46.535 72.965 46.705 ;
        RECT 73.135 46.535 73.425 46.705 ;
        RECT 73.595 46.535 73.885 46.705 ;
        RECT 74.055 46.535 74.345 46.705 ;
        RECT 74.515 46.535 74.805 46.705 ;
        RECT 74.975 46.535 75.265 46.705 ;
        RECT 75.435 46.535 75.725 46.705 ;
        RECT 75.895 46.535 76.185 46.705 ;
        RECT 76.355 46.535 76.645 46.705 ;
        RECT 76.815 46.535 77.105 46.705 ;
        RECT 77.275 46.535 77.565 46.705 ;
        RECT 77.735 46.535 78.025 46.705 ;
        RECT 78.195 46.535 78.485 46.705 ;
        RECT 78.655 46.535 78.945 46.705 ;
        RECT 79.115 46.535 79.405 46.705 ;
        RECT 79.575 46.535 79.865 46.705 ;
        RECT 80.035 46.535 80.325 46.705 ;
        RECT 80.495 46.535 80.785 46.705 ;
        RECT 80.955 46.535 81.245 46.705 ;
        RECT 81.415 46.535 81.705 46.705 ;
        RECT 81.875 46.535 82.165 46.705 ;
        RECT 82.335 46.535 82.625 46.705 ;
        RECT 82.795 46.535 83.085 46.705 ;
        RECT 83.255 46.535 83.545 46.705 ;
        RECT 83.715 46.535 84.005 46.705 ;
        RECT 84.175 46.535 84.465 46.705 ;
        RECT 84.635 46.535 84.925 46.705 ;
        RECT 85.095 46.535 85.385 46.705 ;
        RECT 85.555 46.535 85.845 46.705 ;
        RECT 86.015 46.535 86.305 46.705 ;
        RECT 86.475 46.535 86.765 46.705 ;
        RECT 86.935 46.535 87.225 46.705 ;
        RECT 87.395 46.535 87.685 46.705 ;
        RECT 87.855 46.535 88.145 46.705 ;
        RECT 88.315 46.535 88.605 46.705 ;
        RECT 88.775 46.535 89.065 46.705 ;
        RECT 89.235 46.535 89.525 46.705 ;
        RECT 89.695 46.535 89.985 46.705 ;
        RECT 90.155 46.535 90.445 46.705 ;
        RECT 90.615 46.535 90.905 46.705 ;
        RECT 91.075 46.535 91.365 46.705 ;
        RECT 91.535 46.535 91.825 46.705 ;
        RECT 91.995 46.535 92.285 46.705 ;
        RECT 92.455 46.535 92.745 46.705 ;
        RECT 92.915 46.535 93.205 46.705 ;
        RECT 93.375 46.535 93.665 46.705 ;
        RECT 93.835 46.535 94.125 46.705 ;
        RECT 94.295 46.535 94.585 46.705 ;
        RECT 94.755 46.535 95.045 46.705 ;
        RECT 95.215 46.535 95.505 46.705 ;
        RECT 95.675 46.535 95.965 46.705 ;
        RECT 96.135 46.535 96.425 46.705 ;
        RECT 96.595 46.535 96.885 46.705 ;
        RECT 97.055 46.535 97.345 46.705 ;
        RECT 97.515 46.535 97.805 46.705 ;
        RECT 97.975 46.535 98.265 46.705 ;
        RECT 98.435 46.535 98.725 46.705 ;
        RECT 98.895 46.535 99.185 46.705 ;
        RECT 99.355 46.535 99.645 46.705 ;
        RECT 99.815 46.535 99.960 46.705 ;
        RECT 16.785 45.785 17.995 46.535 ;
        RECT 16.785 45.245 17.305 45.785 ;
        RECT 18.165 45.765 23.510 46.535 ;
        RECT 23.685 45.765 29.030 46.535 ;
        RECT 29.205 45.765 30.875 46.535 ;
        RECT 31.045 45.810 31.335 46.535 ;
        RECT 31.505 45.765 36.850 46.535 ;
        RECT 37.025 45.765 42.370 46.535 ;
        RECT 42.545 45.765 47.890 46.535 ;
        RECT 48.065 45.765 53.410 46.535 ;
        RECT 53.585 45.765 58.930 46.535 ;
        RECT 59.105 45.810 59.395 46.535 ;
        RECT 59.575 46.005 59.905 46.365 ;
        RECT 60.435 46.175 60.765 46.535 ;
        RECT 61.370 46.175 61.700 46.535 ;
      LAYER li1 ;
        RECT 61.010 46.005 61.200 46.105 ;
        RECT 61.870 46.005 62.060 46.365 ;
      LAYER li1 ;
        RECT 62.230 46.175 62.560 46.535 ;
        RECT 59.575 45.815 60.840 46.005 ;
        RECT 17.475 45.075 17.995 45.615 ;
        RECT 18.165 45.245 20.745 45.765 ;
        RECT 20.915 45.075 23.510 45.595 ;
        RECT 23.685 45.245 26.265 45.765 ;
        RECT 26.435 45.075 29.030 45.595 ;
        RECT 29.205 45.245 29.955 45.765 ;
        RECT 30.125 45.075 30.875 45.595 ;
        RECT 31.505 45.245 34.085 45.765 ;
        RECT 16.785 43.985 17.995 45.075 ;
        RECT 18.165 43.985 23.510 45.075 ;
        RECT 23.685 43.985 29.030 45.075 ;
        RECT 29.205 43.985 30.875 45.075 ;
        RECT 31.045 43.985 31.335 45.150 ;
        RECT 34.255 45.075 36.850 45.595 ;
        RECT 37.025 45.245 39.605 45.765 ;
        RECT 39.775 45.075 42.370 45.595 ;
        RECT 42.545 45.245 45.125 45.765 ;
        RECT 45.295 45.075 47.890 45.595 ;
        RECT 48.065 45.245 50.645 45.765 ;
        RECT 50.815 45.075 53.410 45.595 ;
        RECT 53.585 45.245 56.165 45.765 ;
        RECT 56.335 45.075 58.930 45.595 ;
        RECT 31.505 43.985 36.850 45.075 ;
        RECT 37.025 43.985 42.370 45.075 ;
        RECT 42.545 43.985 47.890 45.075 ;
        RECT 48.065 43.985 53.410 45.075 ;
        RECT 53.585 43.985 58.930 45.075 ;
        RECT 59.105 43.985 59.395 45.150 ;
      LAYER li1 ;
        RECT 59.605 45.005 59.915 45.625 ;
      LAYER li1 ;
        RECT 60.630 45.600 60.840 45.815 ;
      LAYER li1 ;
        RECT 61.010 45.775 62.615 46.005 ;
      LAYER li1 ;
        RECT 60.630 45.265 62.165 45.600 ;
        RECT 60.630 45.040 60.840 45.265 ;
      LAYER li1 ;
        RECT 62.335 45.085 62.615 45.775 ;
      LAYER li1 ;
        RECT 62.785 45.765 68.130 46.535 ;
        RECT 68.305 45.765 73.650 46.535 ;
        RECT 73.825 45.765 79.170 46.535 ;
        RECT 79.345 45.765 84.690 46.535 ;
        RECT 84.865 45.765 86.535 46.535 ;
        RECT 87.165 45.810 87.455 46.535 ;
        RECT 87.625 45.765 92.970 46.535 ;
        RECT 93.145 45.765 98.490 46.535 ;
        RECT 98.665 45.785 99.875 46.535 ;
        RECT 62.785 45.245 65.365 45.765 ;
        RECT 60.085 44.870 60.840 45.040 ;
        RECT 59.575 43.985 59.905 44.740 ;
        RECT 60.085 44.155 60.265 44.870 ;
      LAYER li1 ;
        RECT 61.010 44.860 62.615 45.085 ;
      LAYER li1 ;
        RECT 65.535 45.075 68.130 45.595 ;
        RECT 68.305 45.245 70.885 45.765 ;
        RECT 71.055 45.075 73.650 45.595 ;
        RECT 73.825 45.245 76.405 45.765 ;
        RECT 76.575 45.075 79.170 45.595 ;
        RECT 79.345 45.245 81.925 45.765 ;
        RECT 82.095 45.075 84.690 45.595 ;
        RECT 84.865 45.245 85.615 45.765 ;
        RECT 85.785 45.075 86.535 45.595 ;
        RECT 87.625 45.245 90.205 45.765 ;
        RECT 60.470 43.985 60.800 44.685 ;
      LAYER li1 ;
        RECT 61.010 44.155 61.200 44.860 ;
        RECT 61.870 44.855 62.615 44.860 ;
      LAYER li1 ;
        RECT 61.370 43.985 61.700 44.685 ;
      LAYER li1 ;
        RECT 61.870 44.155 62.060 44.855 ;
      LAYER li1 ;
        RECT 62.230 43.985 62.560 44.685 ;
        RECT 62.785 43.985 68.130 45.075 ;
        RECT 68.305 43.985 73.650 45.075 ;
        RECT 73.825 43.985 79.170 45.075 ;
        RECT 79.345 43.985 84.690 45.075 ;
        RECT 84.865 43.985 86.535 45.075 ;
        RECT 87.165 43.985 87.455 45.150 ;
        RECT 90.375 45.075 92.970 45.595 ;
        RECT 93.145 45.245 95.725 45.765 ;
        RECT 95.895 45.075 98.490 45.595 ;
        RECT 87.625 43.985 92.970 45.075 ;
        RECT 93.145 43.985 98.490 45.075 ;
        RECT 98.665 45.075 99.185 45.615 ;
        RECT 99.355 45.245 99.875 45.785 ;
        RECT 98.665 43.985 99.875 45.075 ;
        RECT 16.700 43.815 16.845 43.985 ;
        RECT 17.015 43.815 17.305 43.985 ;
        RECT 17.475 43.815 17.765 43.985 ;
        RECT 17.935 43.815 18.225 43.985 ;
        RECT 18.395 43.815 18.685 43.985 ;
        RECT 18.855 43.815 19.145 43.985 ;
        RECT 19.315 43.815 19.605 43.985 ;
        RECT 19.775 43.815 20.065 43.985 ;
        RECT 20.235 43.815 20.525 43.985 ;
        RECT 20.695 43.815 20.985 43.985 ;
        RECT 21.155 43.815 21.445 43.985 ;
        RECT 21.615 43.815 21.905 43.985 ;
        RECT 22.075 43.815 22.365 43.985 ;
        RECT 22.535 43.815 22.825 43.985 ;
        RECT 22.995 43.815 23.285 43.985 ;
        RECT 23.455 43.815 23.745 43.985 ;
        RECT 23.915 43.815 24.205 43.985 ;
        RECT 24.375 43.815 24.665 43.985 ;
        RECT 24.835 43.815 25.125 43.985 ;
        RECT 25.295 43.815 25.585 43.985 ;
        RECT 25.755 43.815 26.045 43.985 ;
        RECT 26.215 43.815 26.505 43.985 ;
        RECT 26.675 43.815 26.965 43.985 ;
        RECT 27.135 43.815 27.425 43.985 ;
        RECT 27.595 43.815 27.885 43.985 ;
        RECT 28.055 43.815 28.345 43.985 ;
        RECT 28.515 43.815 28.805 43.985 ;
        RECT 28.975 43.815 29.265 43.985 ;
        RECT 29.435 43.815 29.725 43.985 ;
        RECT 29.895 43.815 30.185 43.985 ;
        RECT 30.355 43.815 30.645 43.985 ;
        RECT 30.815 43.815 31.105 43.985 ;
        RECT 31.275 43.815 31.565 43.985 ;
        RECT 31.735 43.815 32.025 43.985 ;
        RECT 32.195 43.815 32.485 43.985 ;
        RECT 32.655 43.815 32.945 43.985 ;
        RECT 33.115 43.815 33.405 43.985 ;
        RECT 33.575 43.815 33.865 43.985 ;
        RECT 34.035 43.815 34.325 43.985 ;
        RECT 34.495 43.815 34.785 43.985 ;
        RECT 34.955 43.815 35.245 43.985 ;
        RECT 35.415 43.815 35.705 43.985 ;
        RECT 35.875 43.815 36.165 43.985 ;
        RECT 36.335 43.815 36.625 43.985 ;
        RECT 36.795 43.815 37.085 43.985 ;
        RECT 37.255 43.815 37.545 43.985 ;
        RECT 37.715 43.815 38.005 43.985 ;
        RECT 38.175 43.815 38.465 43.985 ;
        RECT 38.635 43.815 38.925 43.985 ;
        RECT 39.095 43.815 39.385 43.985 ;
        RECT 39.555 43.815 39.845 43.985 ;
        RECT 40.015 43.815 40.305 43.985 ;
        RECT 40.475 43.815 40.765 43.985 ;
        RECT 40.935 43.815 41.225 43.985 ;
        RECT 41.395 43.815 41.685 43.985 ;
        RECT 41.855 43.815 42.145 43.985 ;
        RECT 42.315 43.815 42.605 43.985 ;
        RECT 42.775 43.815 43.065 43.985 ;
        RECT 43.235 43.815 43.525 43.985 ;
        RECT 43.695 43.815 43.985 43.985 ;
        RECT 44.155 43.815 44.445 43.985 ;
        RECT 44.615 43.815 44.905 43.985 ;
        RECT 45.075 43.815 45.365 43.985 ;
        RECT 45.535 43.815 45.825 43.985 ;
        RECT 45.995 43.815 46.285 43.985 ;
        RECT 46.455 43.815 46.745 43.985 ;
        RECT 46.915 43.815 47.205 43.985 ;
        RECT 47.375 43.815 47.665 43.985 ;
        RECT 47.835 43.815 48.125 43.985 ;
        RECT 48.295 43.815 48.585 43.985 ;
        RECT 48.755 43.815 49.045 43.985 ;
        RECT 49.215 43.815 49.505 43.985 ;
        RECT 49.675 43.815 49.965 43.985 ;
        RECT 50.135 43.815 50.425 43.985 ;
        RECT 50.595 43.815 50.885 43.985 ;
        RECT 51.055 43.815 51.345 43.985 ;
        RECT 51.515 43.815 51.805 43.985 ;
        RECT 51.975 43.815 52.265 43.985 ;
        RECT 52.435 43.815 52.725 43.985 ;
        RECT 52.895 43.815 53.185 43.985 ;
        RECT 53.355 43.815 53.645 43.985 ;
        RECT 53.815 43.815 54.105 43.985 ;
        RECT 54.275 43.815 54.565 43.985 ;
        RECT 54.735 43.815 55.025 43.985 ;
        RECT 55.195 43.815 55.485 43.985 ;
        RECT 55.655 43.815 55.945 43.985 ;
        RECT 56.115 43.815 56.405 43.985 ;
        RECT 56.575 43.815 56.865 43.985 ;
        RECT 57.035 43.815 57.325 43.985 ;
        RECT 57.495 43.815 57.785 43.985 ;
        RECT 57.955 43.815 58.245 43.985 ;
        RECT 58.415 43.815 58.705 43.985 ;
        RECT 58.875 43.815 59.165 43.985 ;
        RECT 59.335 43.815 59.625 43.985 ;
        RECT 59.795 43.815 60.085 43.985 ;
        RECT 60.255 43.815 60.545 43.985 ;
        RECT 60.715 43.815 61.005 43.985 ;
        RECT 61.175 43.815 61.465 43.985 ;
        RECT 61.635 43.815 61.925 43.985 ;
        RECT 62.095 43.815 62.385 43.985 ;
        RECT 62.555 43.815 62.845 43.985 ;
        RECT 63.015 43.815 63.305 43.985 ;
        RECT 63.475 43.815 63.765 43.985 ;
        RECT 63.935 43.815 64.225 43.985 ;
        RECT 64.395 43.815 64.685 43.985 ;
        RECT 64.855 43.815 65.145 43.985 ;
        RECT 65.315 43.815 65.605 43.985 ;
        RECT 65.775 43.815 66.065 43.985 ;
        RECT 66.235 43.815 66.525 43.985 ;
        RECT 66.695 43.815 66.985 43.985 ;
        RECT 67.155 43.815 67.445 43.985 ;
        RECT 67.615 43.815 67.905 43.985 ;
        RECT 68.075 43.815 68.365 43.985 ;
        RECT 68.535 43.815 68.825 43.985 ;
        RECT 68.995 43.815 69.285 43.985 ;
        RECT 69.455 43.815 69.745 43.985 ;
        RECT 69.915 43.815 70.205 43.985 ;
        RECT 70.375 43.815 70.665 43.985 ;
        RECT 70.835 43.815 71.125 43.985 ;
        RECT 71.295 43.815 71.585 43.985 ;
        RECT 71.755 43.815 72.045 43.985 ;
        RECT 72.215 43.815 72.505 43.985 ;
        RECT 72.675 43.815 72.965 43.985 ;
        RECT 73.135 43.815 73.425 43.985 ;
        RECT 73.595 43.815 73.885 43.985 ;
        RECT 74.055 43.815 74.345 43.985 ;
        RECT 74.515 43.815 74.805 43.985 ;
        RECT 74.975 43.815 75.265 43.985 ;
        RECT 75.435 43.815 75.725 43.985 ;
        RECT 75.895 43.815 76.185 43.985 ;
        RECT 76.355 43.815 76.645 43.985 ;
        RECT 76.815 43.815 77.105 43.985 ;
        RECT 77.275 43.815 77.565 43.985 ;
        RECT 77.735 43.815 78.025 43.985 ;
        RECT 78.195 43.815 78.485 43.985 ;
        RECT 78.655 43.815 78.945 43.985 ;
        RECT 79.115 43.815 79.405 43.985 ;
        RECT 79.575 43.815 79.865 43.985 ;
        RECT 80.035 43.815 80.325 43.985 ;
        RECT 80.495 43.815 80.785 43.985 ;
        RECT 80.955 43.815 81.245 43.985 ;
        RECT 81.415 43.815 81.705 43.985 ;
        RECT 81.875 43.815 82.165 43.985 ;
        RECT 82.335 43.815 82.625 43.985 ;
        RECT 82.795 43.815 83.085 43.985 ;
        RECT 83.255 43.815 83.545 43.985 ;
        RECT 83.715 43.815 84.005 43.985 ;
        RECT 84.175 43.815 84.465 43.985 ;
        RECT 84.635 43.815 84.925 43.985 ;
        RECT 85.095 43.815 85.385 43.985 ;
        RECT 85.555 43.815 85.845 43.985 ;
        RECT 86.015 43.815 86.305 43.985 ;
        RECT 86.475 43.815 86.765 43.985 ;
        RECT 86.935 43.815 87.225 43.985 ;
        RECT 87.395 43.815 87.685 43.985 ;
        RECT 87.855 43.815 88.145 43.985 ;
        RECT 88.315 43.815 88.605 43.985 ;
        RECT 88.775 43.815 89.065 43.985 ;
        RECT 89.235 43.815 89.525 43.985 ;
        RECT 89.695 43.815 89.985 43.985 ;
        RECT 90.155 43.815 90.445 43.985 ;
        RECT 90.615 43.815 90.905 43.985 ;
        RECT 91.075 43.815 91.365 43.985 ;
        RECT 91.535 43.815 91.825 43.985 ;
        RECT 91.995 43.815 92.285 43.985 ;
        RECT 92.455 43.815 92.745 43.985 ;
        RECT 92.915 43.815 93.205 43.985 ;
        RECT 93.375 43.815 93.665 43.985 ;
        RECT 93.835 43.815 94.125 43.985 ;
        RECT 94.295 43.815 94.585 43.985 ;
        RECT 94.755 43.815 95.045 43.985 ;
        RECT 95.215 43.815 95.505 43.985 ;
        RECT 95.675 43.815 95.965 43.985 ;
        RECT 96.135 43.815 96.425 43.985 ;
        RECT 96.595 43.815 96.885 43.985 ;
        RECT 97.055 43.815 97.345 43.985 ;
        RECT 97.515 43.815 97.805 43.985 ;
        RECT 97.975 43.815 98.265 43.985 ;
        RECT 98.435 43.815 98.725 43.985 ;
        RECT 98.895 43.815 99.185 43.985 ;
        RECT 99.355 43.815 99.645 43.985 ;
        RECT 99.815 43.815 99.960 43.985 ;
        RECT 16.785 42.725 17.995 43.815 ;
        RECT 18.165 42.725 23.510 43.815 ;
        RECT 23.685 42.725 29.030 43.815 ;
        RECT 29.205 42.725 34.550 43.815 ;
        RECT 34.725 42.725 40.070 43.815 ;
        RECT 40.245 42.725 43.755 43.815 ;
        RECT 16.785 42.015 17.305 42.555 ;
        RECT 17.475 42.185 17.995 42.725 ;
        RECT 18.165 42.035 20.745 42.555 ;
        RECT 20.915 42.205 23.510 42.725 ;
        RECT 23.685 42.035 26.265 42.555 ;
        RECT 26.435 42.205 29.030 42.725 ;
        RECT 29.205 42.035 31.785 42.555 ;
        RECT 31.955 42.205 34.550 42.725 ;
        RECT 34.725 42.035 37.305 42.555 ;
        RECT 37.475 42.205 40.070 42.725 ;
        RECT 40.245 42.035 41.895 42.555 ;
        RECT 42.065 42.205 43.755 42.725 ;
        RECT 44.845 42.650 45.135 43.815 ;
        RECT 45.305 42.725 50.650 43.815 ;
        RECT 50.825 42.725 56.170 43.815 ;
        RECT 56.345 42.725 61.690 43.815 ;
        RECT 61.865 42.725 67.210 43.815 ;
        RECT 67.385 42.725 72.730 43.815 ;
        RECT 45.305 42.035 47.885 42.555 ;
        RECT 48.055 42.205 50.650 42.725 ;
        RECT 50.825 42.035 53.405 42.555 ;
        RECT 53.575 42.205 56.170 42.725 ;
        RECT 56.345 42.035 58.925 42.555 ;
        RECT 59.095 42.205 61.690 42.725 ;
        RECT 61.865 42.035 64.445 42.555 ;
        RECT 64.615 42.205 67.210 42.725 ;
        RECT 67.385 42.035 69.965 42.555 ;
        RECT 70.135 42.205 72.730 42.725 ;
        RECT 72.905 42.650 73.195 43.815 ;
        RECT 73.365 42.725 78.710 43.815 ;
        RECT 78.885 42.725 84.230 43.815 ;
        RECT 84.405 42.725 89.750 43.815 ;
        RECT 89.925 42.725 95.270 43.815 ;
        RECT 95.445 42.725 98.035 43.815 ;
        RECT 73.365 42.035 75.945 42.555 ;
        RECT 76.115 42.205 78.710 42.725 ;
        RECT 78.885 42.035 81.465 42.555 ;
        RECT 81.635 42.205 84.230 42.725 ;
        RECT 84.405 42.035 86.985 42.555 ;
        RECT 87.155 42.205 89.750 42.725 ;
        RECT 89.925 42.035 92.505 42.555 ;
        RECT 92.675 42.205 95.270 42.725 ;
        RECT 95.445 42.035 96.655 42.555 ;
        RECT 96.825 42.205 98.035 42.725 ;
        RECT 98.665 42.725 99.875 43.815 ;
        RECT 98.665 42.185 99.185 42.725 ;
        RECT 16.785 41.265 17.995 42.015 ;
        RECT 18.165 41.265 23.510 42.035 ;
        RECT 23.685 41.265 29.030 42.035 ;
        RECT 29.205 41.265 34.550 42.035 ;
        RECT 34.725 41.265 40.070 42.035 ;
        RECT 40.245 41.265 43.755 42.035 ;
        RECT 44.845 41.265 45.135 41.990 ;
        RECT 45.305 41.265 50.650 42.035 ;
        RECT 50.825 41.265 56.170 42.035 ;
        RECT 56.345 41.265 61.690 42.035 ;
        RECT 61.865 41.265 67.210 42.035 ;
        RECT 67.385 41.265 72.730 42.035 ;
        RECT 72.905 41.265 73.195 41.990 ;
        RECT 73.365 41.265 78.710 42.035 ;
        RECT 78.885 41.265 84.230 42.035 ;
        RECT 84.405 41.265 89.750 42.035 ;
        RECT 89.925 41.265 95.270 42.035 ;
        RECT 95.445 41.265 98.035 42.035 ;
        RECT 99.355 42.015 99.875 42.555 ;
        RECT 98.665 41.265 99.875 42.015 ;
        RECT 16.700 41.095 16.845 41.265 ;
        RECT 17.015 41.095 17.305 41.265 ;
        RECT 17.475 41.095 17.765 41.265 ;
        RECT 17.935 41.095 18.225 41.265 ;
        RECT 18.395 41.095 18.685 41.265 ;
        RECT 18.855 41.095 19.145 41.265 ;
        RECT 19.315 41.095 19.605 41.265 ;
        RECT 19.775 41.095 20.065 41.265 ;
        RECT 20.235 41.095 20.525 41.265 ;
        RECT 20.695 41.095 20.985 41.265 ;
        RECT 21.155 41.095 21.445 41.265 ;
        RECT 21.615 41.095 21.905 41.265 ;
        RECT 22.075 41.095 22.365 41.265 ;
        RECT 22.535 41.095 22.825 41.265 ;
        RECT 22.995 41.095 23.285 41.265 ;
        RECT 23.455 41.095 23.745 41.265 ;
        RECT 23.915 41.095 24.205 41.265 ;
        RECT 24.375 41.095 24.665 41.265 ;
        RECT 24.835 41.095 25.125 41.265 ;
        RECT 25.295 41.095 25.585 41.265 ;
        RECT 25.755 41.095 26.045 41.265 ;
        RECT 26.215 41.095 26.505 41.265 ;
        RECT 26.675 41.095 26.965 41.265 ;
        RECT 27.135 41.095 27.425 41.265 ;
        RECT 27.595 41.095 27.885 41.265 ;
        RECT 28.055 41.095 28.345 41.265 ;
        RECT 28.515 41.095 28.805 41.265 ;
        RECT 28.975 41.095 29.265 41.265 ;
        RECT 29.435 41.095 29.725 41.265 ;
        RECT 29.895 41.095 30.185 41.265 ;
        RECT 30.355 41.095 30.645 41.265 ;
        RECT 30.815 41.095 31.105 41.265 ;
        RECT 31.275 41.095 31.565 41.265 ;
        RECT 31.735 41.095 32.025 41.265 ;
        RECT 32.195 41.095 32.485 41.265 ;
        RECT 32.655 41.095 32.945 41.265 ;
        RECT 33.115 41.095 33.405 41.265 ;
        RECT 33.575 41.095 33.865 41.265 ;
        RECT 34.035 41.095 34.325 41.265 ;
        RECT 34.495 41.095 34.785 41.265 ;
        RECT 34.955 41.095 35.245 41.265 ;
        RECT 35.415 41.095 35.705 41.265 ;
        RECT 35.875 41.095 36.165 41.265 ;
        RECT 36.335 41.095 36.625 41.265 ;
        RECT 36.795 41.095 37.085 41.265 ;
        RECT 37.255 41.095 37.545 41.265 ;
        RECT 37.715 41.095 38.005 41.265 ;
        RECT 38.175 41.095 38.465 41.265 ;
        RECT 38.635 41.095 38.925 41.265 ;
        RECT 39.095 41.095 39.385 41.265 ;
        RECT 39.555 41.095 39.845 41.265 ;
        RECT 40.015 41.095 40.305 41.265 ;
        RECT 40.475 41.095 40.765 41.265 ;
        RECT 40.935 41.095 41.225 41.265 ;
        RECT 41.395 41.095 41.685 41.265 ;
        RECT 41.855 41.095 42.145 41.265 ;
        RECT 42.315 41.095 42.605 41.265 ;
        RECT 42.775 41.095 43.065 41.265 ;
        RECT 43.235 41.095 43.525 41.265 ;
        RECT 43.695 41.095 43.985 41.265 ;
        RECT 44.155 41.095 44.445 41.265 ;
        RECT 44.615 41.095 44.905 41.265 ;
        RECT 45.075 41.095 45.365 41.265 ;
        RECT 45.535 41.095 45.825 41.265 ;
        RECT 45.995 41.095 46.285 41.265 ;
        RECT 46.455 41.095 46.745 41.265 ;
        RECT 46.915 41.095 47.205 41.265 ;
        RECT 47.375 41.095 47.665 41.265 ;
        RECT 47.835 41.095 48.125 41.265 ;
        RECT 48.295 41.095 48.585 41.265 ;
        RECT 48.755 41.095 49.045 41.265 ;
        RECT 49.215 41.095 49.505 41.265 ;
        RECT 49.675 41.095 49.965 41.265 ;
        RECT 50.135 41.095 50.425 41.265 ;
        RECT 50.595 41.095 50.885 41.265 ;
        RECT 51.055 41.095 51.345 41.265 ;
        RECT 51.515 41.095 51.805 41.265 ;
        RECT 51.975 41.095 52.265 41.265 ;
        RECT 52.435 41.095 52.725 41.265 ;
        RECT 52.895 41.095 53.185 41.265 ;
        RECT 53.355 41.095 53.645 41.265 ;
        RECT 53.815 41.095 54.105 41.265 ;
        RECT 54.275 41.095 54.565 41.265 ;
        RECT 54.735 41.095 55.025 41.265 ;
        RECT 55.195 41.095 55.485 41.265 ;
        RECT 55.655 41.095 55.945 41.265 ;
        RECT 56.115 41.095 56.405 41.265 ;
        RECT 56.575 41.095 56.865 41.265 ;
        RECT 57.035 41.095 57.325 41.265 ;
        RECT 57.495 41.095 57.785 41.265 ;
        RECT 57.955 41.095 58.245 41.265 ;
        RECT 58.415 41.095 58.705 41.265 ;
        RECT 58.875 41.095 59.165 41.265 ;
        RECT 59.335 41.095 59.625 41.265 ;
        RECT 59.795 41.095 60.085 41.265 ;
        RECT 60.255 41.095 60.545 41.265 ;
        RECT 60.715 41.095 61.005 41.265 ;
        RECT 61.175 41.095 61.465 41.265 ;
        RECT 61.635 41.095 61.925 41.265 ;
        RECT 62.095 41.095 62.385 41.265 ;
        RECT 62.555 41.095 62.845 41.265 ;
        RECT 63.015 41.095 63.305 41.265 ;
        RECT 63.475 41.095 63.765 41.265 ;
        RECT 63.935 41.095 64.225 41.265 ;
        RECT 64.395 41.095 64.685 41.265 ;
        RECT 64.855 41.095 65.145 41.265 ;
        RECT 65.315 41.095 65.605 41.265 ;
        RECT 65.775 41.095 66.065 41.265 ;
        RECT 66.235 41.095 66.525 41.265 ;
        RECT 66.695 41.095 66.985 41.265 ;
        RECT 67.155 41.095 67.445 41.265 ;
        RECT 67.615 41.095 67.905 41.265 ;
        RECT 68.075 41.095 68.365 41.265 ;
        RECT 68.535 41.095 68.825 41.265 ;
        RECT 68.995 41.095 69.285 41.265 ;
        RECT 69.455 41.095 69.745 41.265 ;
        RECT 69.915 41.095 70.205 41.265 ;
        RECT 70.375 41.095 70.665 41.265 ;
        RECT 70.835 41.095 71.125 41.265 ;
        RECT 71.295 41.095 71.585 41.265 ;
        RECT 71.755 41.095 72.045 41.265 ;
        RECT 72.215 41.095 72.505 41.265 ;
        RECT 72.675 41.095 72.965 41.265 ;
        RECT 73.135 41.095 73.425 41.265 ;
        RECT 73.595 41.095 73.885 41.265 ;
        RECT 74.055 41.095 74.345 41.265 ;
        RECT 74.515 41.095 74.805 41.265 ;
        RECT 74.975 41.095 75.265 41.265 ;
        RECT 75.435 41.095 75.725 41.265 ;
        RECT 75.895 41.095 76.185 41.265 ;
        RECT 76.355 41.095 76.645 41.265 ;
        RECT 76.815 41.095 77.105 41.265 ;
        RECT 77.275 41.095 77.565 41.265 ;
        RECT 77.735 41.095 78.025 41.265 ;
        RECT 78.195 41.095 78.485 41.265 ;
        RECT 78.655 41.095 78.945 41.265 ;
        RECT 79.115 41.095 79.405 41.265 ;
        RECT 79.575 41.095 79.865 41.265 ;
        RECT 80.035 41.095 80.325 41.265 ;
        RECT 80.495 41.095 80.785 41.265 ;
        RECT 80.955 41.095 81.245 41.265 ;
        RECT 81.415 41.095 81.705 41.265 ;
        RECT 81.875 41.095 82.165 41.265 ;
        RECT 82.335 41.095 82.625 41.265 ;
        RECT 82.795 41.095 83.085 41.265 ;
        RECT 83.255 41.095 83.545 41.265 ;
        RECT 83.715 41.095 84.005 41.265 ;
        RECT 84.175 41.095 84.465 41.265 ;
        RECT 84.635 41.095 84.925 41.265 ;
        RECT 85.095 41.095 85.385 41.265 ;
        RECT 85.555 41.095 85.845 41.265 ;
        RECT 86.015 41.095 86.305 41.265 ;
        RECT 86.475 41.095 86.765 41.265 ;
        RECT 86.935 41.095 87.225 41.265 ;
        RECT 87.395 41.095 87.685 41.265 ;
        RECT 87.855 41.095 88.145 41.265 ;
        RECT 88.315 41.095 88.605 41.265 ;
        RECT 88.775 41.095 89.065 41.265 ;
        RECT 89.235 41.095 89.525 41.265 ;
        RECT 89.695 41.095 89.985 41.265 ;
        RECT 90.155 41.095 90.445 41.265 ;
        RECT 90.615 41.095 90.905 41.265 ;
        RECT 91.075 41.095 91.365 41.265 ;
        RECT 91.535 41.095 91.825 41.265 ;
        RECT 91.995 41.095 92.285 41.265 ;
        RECT 92.455 41.095 92.745 41.265 ;
        RECT 92.915 41.095 93.205 41.265 ;
        RECT 93.375 41.095 93.665 41.265 ;
        RECT 93.835 41.095 94.125 41.265 ;
        RECT 94.295 41.095 94.585 41.265 ;
        RECT 94.755 41.095 95.045 41.265 ;
        RECT 95.215 41.095 95.505 41.265 ;
        RECT 95.675 41.095 95.965 41.265 ;
        RECT 96.135 41.095 96.425 41.265 ;
        RECT 96.595 41.095 96.885 41.265 ;
        RECT 97.055 41.095 97.345 41.265 ;
        RECT 97.515 41.095 97.805 41.265 ;
        RECT 97.975 41.095 98.265 41.265 ;
        RECT 98.435 41.095 98.725 41.265 ;
        RECT 98.895 41.095 99.185 41.265 ;
        RECT 99.355 41.095 99.645 41.265 ;
        RECT 99.815 41.095 99.960 41.265 ;
        RECT 16.785 40.345 17.995 41.095 ;
        RECT 16.785 39.805 17.305 40.345 ;
        RECT 18.165 40.325 23.510 41.095 ;
        RECT 23.685 40.325 29.030 41.095 ;
        RECT 29.205 40.325 30.875 41.095 ;
        RECT 31.045 40.370 31.335 41.095 ;
        RECT 31.505 40.325 36.850 41.095 ;
        RECT 37.025 40.325 42.370 41.095 ;
        RECT 42.545 40.325 47.890 41.095 ;
        RECT 48.065 40.325 53.410 41.095 ;
        RECT 53.585 40.325 58.930 41.095 ;
        RECT 59.105 40.370 59.395 41.095 ;
        RECT 59.565 40.325 64.910 41.095 ;
        RECT 65.085 40.325 70.430 41.095 ;
        RECT 70.605 40.325 75.950 41.095 ;
        RECT 76.125 40.325 81.470 41.095 ;
        RECT 81.645 40.325 86.990 41.095 ;
        RECT 87.165 40.370 87.455 41.095 ;
        RECT 87.625 40.325 92.970 41.095 ;
        RECT 93.145 40.325 98.490 41.095 ;
        RECT 98.665 40.345 99.875 41.095 ;
        RECT 17.475 39.635 17.995 40.175 ;
        RECT 18.165 39.805 20.745 40.325 ;
        RECT 20.915 39.635 23.510 40.155 ;
        RECT 23.685 39.805 26.265 40.325 ;
        RECT 26.435 39.635 29.030 40.155 ;
        RECT 29.205 39.805 29.955 40.325 ;
        RECT 30.125 39.635 30.875 40.155 ;
        RECT 31.505 39.805 34.085 40.325 ;
        RECT 16.785 38.545 17.995 39.635 ;
        RECT 18.165 38.545 23.510 39.635 ;
        RECT 23.685 38.545 29.030 39.635 ;
        RECT 29.205 38.545 30.875 39.635 ;
        RECT 31.045 38.545 31.335 39.710 ;
        RECT 34.255 39.635 36.850 40.155 ;
        RECT 37.025 39.805 39.605 40.325 ;
        RECT 39.775 39.635 42.370 40.155 ;
        RECT 42.545 39.805 45.125 40.325 ;
        RECT 45.295 39.635 47.890 40.155 ;
        RECT 48.065 39.805 50.645 40.325 ;
        RECT 50.815 39.635 53.410 40.155 ;
        RECT 53.585 39.805 56.165 40.325 ;
        RECT 56.335 39.635 58.930 40.155 ;
        RECT 59.565 39.805 62.145 40.325 ;
        RECT 31.505 38.545 36.850 39.635 ;
        RECT 37.025 38.545 42.370 39.635 ;
        RECT 42.545 38.545 47.890 39.635 ;
        RECT 48.065 38.545 53.410 39.635 ;
        RECT 53.585 38.545 58.930 39.635 ;
        RECT 59.105 38.545 59.395 39.710 ;
        RECT 62.315 39.635 64.910 40.155 ;
        RECT 65.085 39.805 67.665 40.325 ;
        RECT 67.835 39.635 70.430 40.155 ;
        RECT 70.605 39.805 73.185 40.325 ;
        RECT 73.355 39.635 75.950 40.155 ;
        RECT 76.125 39.805 78.705 40.325 ;
        RECT 78.875 39.635 81.470 40.155 ;
        RECT 81.645 39.805 84.225 40.325 ;
        RECT 84.395 39.635 86.990 40.155 ;
        RECT 87.625 39.805 90.205 40.325 ;
        RECT 59.565 38.545 64.910 39.635 ;
        RECT 65.085 38.545 70.430 39.635 ;
        RECT 70.605 38.545 75.950 39.635 ;
        RECT 76.125 38.545 81.470 39.635 ;
        RECT 81.645 38.545 86.990 39.635 ;
        RECT 87.165 38.545 87.455 39.710 ;
        RECT 90.375 39.635 92.970 40.155 ;
        RECT 93.145 39.805 95.725 40.325 ;
        RECT 95.895 39.635 98.490 40.155 ;
        RECT 87.625 38.545 92.970 39.635 ;
        RECT 93.145 38.545 98.490 39.635 ;
        RECT 98.665 39.635 99.185 40.175 ;
        RECT 99.355 39.805 99.875 40.345 ;
        RECT 98.665 38.545 99.875 39.635 ;
        RECT 16.700 38.375 16.845 38.545 ;
        RECT 17.015 38.375 17.305 38.545 ;
        RECT 17.475 38.375 17.765 38.545 ;
        RECT 17.935 38.375 18.225 38.545 ;
        RECT 18.395 38.375 18.685 38.545 ;
        RECT 18.855 38.375 19.145 38.545 ;
        RECT 19.315 38.375 19.605 38.545 ;
        RECT 19.775 38.375 20.065 38.545 ;
        RECT 20.235 38.375 20.525 38.545 ;
        RECT 20.695 38.375 20.985 38.545 ;
        RECT 21.155 38.375 21.445 38.545 ;
        RECT 21.615 38.375 21.905 38.545 ;
        RECT 22.075 38.375 22.365 38.545 ;
        RECT 22.535 38.375 22.825 38.545 ;
        RECT 22.995 38.375 23.285 38.545 ;
        RECT 23.455 38.375 23.745 38.545 ;
        RECT 23.915 38.375 24.205 38.545 ;
        RECT 24.375 38.375 24.665 38.545 ;
        RECT 24.835 38.375 25.125 38.545 ;
        RECT 25.295 38.375 25.585 38.545 ;
        RECT 25.755 38.375 26.045 38.545 ;
        RECT 26.215 38.375 26.505 38.545 ;
        RECT 26.675 38.375 26.965 38.545 ;
        RECT 27.135 38.375 27.425 38.545 ;
        RECT 27.595 38.375 27.885 38.545 ;
        RECT 28.055 38.375 28.345 38.545 ;
        RECT 28.515 38.375 28.805 38.545 ;
        RECT 28.975 38.375 29.265 38.545 ;
        RECT 29.435 38.375 29.725 38.545 ;
        RECT 29.895 38.375 30.185 38.545 ;
        RECT 30.355 38.375 30.645 38.545 ;
        RECT 30.815 38.375 31.105 38.545 ;
        RECT 31.275 38.375 31.565 38.545 ;
        RECT 31.735 38.375 32.025 38.545 ;
        RECT 32.195 38.375 32.485 38.545 ;
        RECT 32.655 38.375 32.945 38.545 ;
        RECT 33.115 38.375 33.405 38.545 ;
        RECT 33.575 38.375 33.865 38.545 ;
        RECT 34.035 38.375 34.325 38.545 ;
        RECT 34.495 38.375 34.785 38.545 ;
        RECT 34.955 38.375 35.245 38.545 ;
        RECT 35.415 38.375 35.705 38.545 ;
        RECT 35.875 38.375 36.165 38.545 ;
        RECT 36.335 38.375 36.625 38.545 ;
        RECT 36.795 38.375 37.085 38.545 ;
        RECT 37.255 38.375 37.545 38.545 ;
        RECT 37.715 38.375 38.005 38.545 ;
        RECT 38.175 38.375 38.465 38.545 ;
        RECT 38.635 38.375 38.925 38.545 ;
        RECT 39.095 38.375 39.385 38.545 ;
        RECT 39.555 38.375 39.845 38.545 ;
        RECT 40.015 38.375 40.305 38.545 ;
        RECT 40.475 38.375 40.765 38.545 ;
        RECT 40.935 38.375 41.225 38.545 ;
        RECT 41.395 38.375 41.685 38.545 ;
        RECT 41.855 38.375 42.145 38.545 ;
        RECT 42.315 38.375 42.605 38.545 ;
        RECT 42.775 38.375 43.065 38.545 ;
        RECT 43.235 38.375 43.525 38.545 ;
        RECT 43.695 38.375 43.985 38.545 ;
        RECT 44.155 38.375 44.445 38.545 ;
        RECT 44.615 38.375 44.905 38.545 ;
        RECT 45.075 38.375 45.365 38.545 ;
        RECT 45.535 38.375 45.825 38.545 ;
        RECT 45.995 38.375 46.285 38.545 ;
        RECT 46.455 38.375 46.745 38.545 ;
        RECT 46.915 38.375 47.205 38.545 ;
        RECT 47.375 38.375 47.665 38.545 ;
        RECT 47.835 38.375 48.125 38.545 ;
        RECT 48.295 38.375 48.585 38.545 ;
        RECT 48.755 38.375 49.045 38.545 ;
        RECT 49.215 38.375 49.505 38.545 ;
        RECT 49.675 38.375 49.965 38.545 ;
        RECT 50.135 38.375 50.425 38.545 ;
        RECT 50.595 38.375 50.885 38.545 ;
        RECT 51.055 38.375 51.345 38.545 ;
        RECT 51.515 38.375 51.805 38.545 ;
        RECT 51.975 38.375 52.265 38.545 ;
        RECT 52.435 38.375 52.725 38.545 ;
        RECT 52.895 38.375 53.185 38.545 ;
        RECT 53.355 38.375 53.645 38.545 ;
        RECT 53.815 38.375 54.105 38.545 ;
        RECT 54.275 38.375 54.565 38.545 ;
        RECT 54.735 38.375 55.025 38.545 ;
        RECT 55.195 38.375 55.485 38.545 ;
        RECT 55.655 38.375 55.945 38.545 ;
        RECT 56.115 38.375 56.405 38.545 ;
        RECT 56.575 38.375 56.865 38.545 ;
        RECT 57.035 38.375 57.325 38.545 ;
        RECT 57.495 38.375 57.785 38.545 ;
        RECT 57.955 38.375 58.245 38.545 ;
        RECT 58.415 38.375 58.705 38.545 ;
        RECT 58.875 38.375 59.165 38.545 ;
        RECT 59.335 38.375 59.625 38.545 ;
        RECT 59.795 38.375 60.085 38.545 ;
        RECT 60.255 38.375 60.545 38.545 ;
        RECT 60.715 38.375 61.005 38.545 ;
        RECT 61.175 38.375 61.465 38.545 ;
        RECT 61.635 38.375 61.925 38.545 ;
        RECT 62.095 38.375 62.385 38.545 ;
        RECT 62.555 38.375 62.845 38.545 ;
        RECT 63.015 38.375 63.305 38.545 ;
        RECT 63.475 38.375 63.765 38.545 ;
        RECT 63.935 38.375 64.225 38.545 ;
        RECT 64.395 38.375 64.685 38.545 ;
        RECT 64.855 38.375 65.145 38.545 ;
        RECT 65.315 38.375 65.605 38.545 ;
        RECT 65.775 38.375 66.065 38.545 ;
        RECT 66.235 38.375 66.525 38.545 ;
        RECT 66.695 38.375 66.985 38.545 ;
        RECT 67.155 38.375 67.445 38.545 ;
        RECT 67.615 38.375 67.905 38.545 ;
        RECT 68.075 38.375 68.365 38.545 ;
        RECT 68.535 38.375 68.825 38.545 ;
        RECT 68.995 38.375 69.285 38.545 ;
        RECT 69.455 38.375 69.745 38.545 ;
        RECT 69.915 38.375 70.205 38.545 ;
        RECT 70.375 38.375 70.665 38.545 ;
        RECT 70.835 38.375 71.125 38.545 ;
        RECT 71.295 38.375 71.585 38.545 ;
        RECT 71.755 38.375 72.045 38.545 ;
        RECT 72.215 38.375 72.505 38.545 ;
        RECT 72.675 38.375 72.965 38.545 ;
        RECT 73.135 38.375 73.425 38.545 ;
        RECT 73.595 38.375 73.885 38.545 ;
        RECT 74.055 38.375 74.345 38.545 ;
        RECT 74.515 38.375 74.805 38.545 ;
        RECT 74.975 38.375 75.265 38.545 ;
        RECT 75.435 38.375 75.725 38.545 ;
        RECT 75.895 38.375 76.185 38.545 ;
        RECT 76.355 38.375 76.645 38.545 ;
        RECT 76.815 38.375 77.105 38.545 ;
        RECT 77.275 38.375 77.565 38.545 ;
        RECT 77.735 38.375 78.025 38.545 ;
        RECT 78.195 38.375 78.485 38.545 ;
        RECT 78.655 38.375 78.945 38.545 ;
        RECT 79.115 38.375 79.405 38.545 ;
        RECT 79.575 38.375 79.865 38.545 ;
        RECT 80.035 38.375 80.325 38.545 ;
        RECT 80.495 38.375 80.785 38.545 ;
        RECT 80.955 38.375 81.245 38.545 ;
        RECT 81.415 38.375 81.705 38.545 ;
        RECT 81.875 38.375 82.165 38.545 ;
        RECT 82.335 38.375 82.625 38.545 ;
        RECT 82.795 38.375 83.085 38.545 ;
        RECT 83.255 38.375 83.545 38.545 ;
        RECT 83.715 38.375 84.005 38.545 ;
        RECT 84.175 38.375 84.465 38.545 ;
        RECT 84.635 38.375 84.925 38.545 ;
        RECT 85.095 38.375 85.385 38.545 ;
        RECT 85.555 38.375 85.845 38.545 ;
        RECT 86.015 38.375 86.305 38.545 ;
        RECT 86.475 38.375 86.765 38.545 ;
        RECT 86.935 38.375 87.225 38.545 ;
        RECT 87.395 38.375 87.685 38.545 ;
        RECT 87.855 38.375 88.145 38.545 ;
        RECT 88.315 38.375 88.605 38.545 ;
        RECT 88.775 38.375 89.065 38.545 ;
        RECT 89.235 38.375 89.525 38.545 ;
        RECT 89.695 38.375 89.985 38.545 ;
        RECT 90.155 38.375 90.445 38.545 ;
        RECT 90.615 38.375 90.905 38.545 ;
        RECT 91.075 38.375 91.365 38.545 ;
        RECT 91.535 38.375 91.825 38.545 ;
        RECT 91.995 38.375 92.285 38.545 ;
        RECT 92.455 38.375 92.745 38.545 ;
        RECT 92.915 38.375 93.205 38.545 ;
        RECT 93.375 38.375 93.665 38.545 ;
        RECT 93.835 38.375 94.125 38.545 ;
        RECT 94.295 38.375 94.585 38.545 ;
        RECT 94.755 38.375 95.045 38.545 ;
        RECT 95.215 38.375 95.505 38.545 ;
        RECT 95.675 38.375 95.965 38.545 ;
        RECT 96.135 38.375 96.425 38.545 ;
        RECT 96.595 38.375 96.885 38.545 ;
        RECT 97.055 38.375 97.345 38.545 ;
        RECT 97.515 38.375 97.805 38.545 ;
        RECT 97.975 38.375 98.265 38.545 ;
        RECT 98.435 38.375 98.725 38.545 ;
        RECT 98.895 38.375 99.185 38.545 ;
        RECT 99.355 38.375 99.645 38.545 ;
        RECT 99.815 38.375 99.960 38.545 ;
        RECT 16.785 37.285 17.995 38.375 ;
        RECT 18.165 37.285 23.510 38.375 ;
        RECT 23.685 37.285 29.030 38.375 ;
        RECT 29.205 37.285 34.550 38.375 ;
        RECT 34.725 37.285 40.070 38.375 ;
        RECT 40.245 37.285 43.755 38.375 ;
        RECT 16.785 36.575 17.305 37.115 ;
        RECT 17.475 36.745 17.995 37.285 ;
        RECT 18.165 36.595 20.745 37.115 ;
        RECT 20.915 36.765 23.510 37.285 ;
        RECT 23.685 36.595 26.265 37.115 ;
        RECT 26.435 36.765 29.030 37.285 ;
        RECT 29.205 36.595 31.785 37.115 ;
        RECT 31.955 36.765 34.550 37.285 ;
        RECT 34.725 36.595 37.305 37.115 ;
        RECT 37.475 36.765 40.070 37.285 ;
        RECT 40.245 36.595 41.895 37.115 ;
        RECT 42.065 36.765 43.755 37.285 ;
        RECT 44.845 37.210 45.135 38.375 ;
        RECT 45.305 37.285 50.650 38.375 ;
        RECT 50.825 37.285 56.170 38.375 ;
        RECT 56.345 37.285 61.690 38.375 ;
        RECT 61.865 37.285 67.210 38.375 ;
        RECT 67.385 37.285 72.730 38.375 ;
        RECT 45.305 36.595 47.885 37.115 ;
        RECT 48.055 36.765 50.650 37.285 ;
        RECT 50.825 36.595 53.405 37.115 ;
        RECT 53.575 36.765 56.170 37.285 ;
        RECT 56.345 36.595 58.925 37.115 ;
        RECT 59.095 36.765 61.690 37.285 ;
        RECT 61.865 36.595 64.445 37.115 ;
        RECT 64.615 36.765 67.210 37.285 ;
        RECT 67.385 36.595 69.965 37.115 ;
        RECT 70.135 36.765 72.730 37.285 ;
        RECT 72.905 37.210 73.195 38.375 ;
        RECT 73.365 37.285 78.710 38.375 ;
        RECT 78.885 37.285 84.230 38.375 ;
        RECT 84.405 37.285 89.750 38.375 ;
        RECT 89.925 37.285 93.435 38.375 ;
        RECT 93.795 37.650 94.125 38.375 ;
        RECT 73.365 36.595 75.945 37.115 ;
        RECT 76.115 36.765 78.710 37.285 ;
        RECT 78.885 36.595 81.465 37.115 ;
        RECT 81.635 36.765 84.230 37.285 ;
        RECT 84.405 36.595 86.985 37.115 ;
        RECT 87.155 36.765 89.750 37.285 ;
        RECT 89.925 36.595 91.575 37.115 ;
        RECT 91.745 36.765 93.435 37.285 ;
        RECT 16.785 35.825 17.995 36.575 ;
        RECT 18.165 35.825 23.510 36.595 ;
        RECT 23.685 35.825 29.030 36.595 ;
        RECT 29.205 35.825 34.550 36.595 ;
        RECT 34.725 35.825 40.070 36.595 ;
        RECT 40.245 35.825 43.755 36.595 ;
        RECT 44.845 35.825 45.135 36.550 ;
        RECT 45.305 35.825 50.650 36.595 ;
        RECT 50.825 35.825 56.170 36.595 ;
        RECT 56.345 35.825 61.690 36.595 ;
        RECT 61.865 35.825 67.210 36.595 ;
        RECT 67.385 35.825 72.730 36.595 ;
        RECT 72.905 35.825 73.195 36.550 ;
        RECT 73.365 35.825 78.710 36.595 ;
        RECT 78.885 35.825 84.230 36.595 ;
        RECT 84.405 35.825 89.750 36.595 ;
        RECT 89.925 35.825 93.435 36.595 ;
      LAYER li1 ;
        RECT 93.605 35.995 94.125 37.480 ;
      LAYER li1 ;
        RECT 94.985 37.285 98.495 38.375 ;
        RECT 94.985 36.595 96.635 37.115 ;
        RECT 96.805 36.765 98.495 37.285 ;
        RECT 98.665 37.285 99.875 38.375 ;
        RECT 98.665 36.745 99.185 37.285 ;
        RECT 94.295 35.825 94.635 36.485 ;
        RECT 94.985 35.825 98.495 36.595 ;
        RECT 99.355 36.575 99.875 37.115 ;
        RECT 98.665 35.825 99.875 36.575 ;
        RECT 16.700 35.655 16.845 35.825 ;
        RECT 17.015 35.655 17.305 35.825 ;
        RECT 17.475 35.655 17.765 35.825 ;
        RECT 17.935 35.655 18.225 35.825 ;
        RECT 18.395 35.655 18.685 35.825 ;
        RECT 18.855 35.655 19.145 35.825 ;
        RECT 19.315 35.655 19.605 35.825 ;
        RECT 19.775 35.655 20.065 35.825 ;
        RECT 20.235 35.655 20.525 35.825 ;
        RECT 20.695 35.655 20.985 35.825 ;
        RECT 21.155 35.655 21.445 35.825 ;
        RECT 21.615 35.655 21.905 35.825 ;
        RECT 22.075 35.655 22.365 35.825 ;
        RECT 22.535 35.655 22.825 35.825 ;
        RECT 22.995 35.655 23.285 35.825 ;
        RECT 23.455 35.655 23.745 35.825 ;
        RECT 23.915 35.655 24.205 35.825 ;
        RECT 24.375 35.655 24.665 35.825 ;
        RECT 24.835 35.655 25.125 35.825 ;
        RECT 25.295 35.655 25.585 35.825 ;
        RECT 25.755 35.655 26.045 35.825 ;
        RECT 26.215 35.655 26.505 35.825 ;
        RECT 26.675 35.655 26.965 35.825 ;
        RECT 27.135 35.655 27.425 35.825 ;
        RECT 27.595 35.655 27.885 35.825 ;
        RECT 28.055 35.655 28.345 35.825 ;
        RECT 28.515 35.655 28.805 35.825 ;
        RECT 28.975 35.655 29.265 35.825 ;
        RECT 29.435 35.655 29.725 35.825 ;
        RECT 29.895 35.655 30.185 35.825 ;
        RECT 30.355 35.655 30.645 35.825 ;
        RECT 30.815 35.655 31.105 35.825 ;
        RECT 31.275 35.655 31.565 35.825 ;
        RECT 31.735 35.655 32.025 35.825 ;
        RECT 32.195 35.655 32.485 35.825 ;
        RECT 32.655 35.655 32.945 35.825 ;
        RECT 33.115 35.655 33.405 35.825 ;
        RECT 33.575 35.655 33.865 35.825 ;
        RECT 34.035 35.655 34.325 35.825 ;
        RECT 34.495 35.655 34.785 35.825 ;
        RECT 34.955 35.655 35.245 35.825 ;
        RECT 35.415 35.655 35.705 35.825 ;
        RECT 35.875 35.655 36.165 35.825 ;
        RECT 36.335 35.655 36.625 35.825 ;
        RECT 36.795 35.655 37.085 35.825 ;
        RECT 37.255 35.655 37.545 35.825 ;
        RECT 37.715 35.655 38.005 35.825 ;
        RECT 38.175 35.655 38.465 35.825 ;
        RECT 38.635 35.655 38.925 35.825 ;
        RECT 39.095 35.655 39.385 35.825 ;
        RECT 39.555 35.655 39.845 35.825 ;
        RECT 40.015 35.655 40.305 35.825 ;
        RECT 40.475 35.655 40.765 35.825 ;
        RECT 40.935 35.655 41.225 35.825 ;
        RECT 41.395 35.655 41.685 35.825 ;
        RECT 41.855 35.655 42.145 35.825 ;
        RECT 42.315 35.655 42.605 35.825 ;
        RECT 42.775 35.655 43.065 35.825 ;
        RECT 43.235 35.655 43.525 35.825 ;
        RECT 43.695 35.655 43.985 35.825 ;
        RECT 44.155 35.655 44.445 35.825 ;
        RECT 44.615 35.655 44.905 35.825 ;
        RECT 45.075 35.655 45.365 35.825 ;
        RECT 45.535 35.655 45.825 35.825 ;
        RECT 45.995 35.655 46.285 35.825 ;
        RECT 46.455 35.655 46.745 35.825 ;
        RECT 46.915 35.655 47.205 35.825 ;
        RECT 47.375 35.655 47.665 35.825 ;
        RECT 47.835 35.655 48.125 35.825 ;
        RECT 48.295 35.655 48.585 35.825 ;
        RECT 48.755 35.655 49.045 35.825 ;
        RECT 49.215 35.655 49.505 35.825 ;
        RECT 49.675 35.655 49.965 35.825 ;
        RECT 50.135 35.655 50.425 35.825 ;
        RECT 50.595 35.655 50.885 35.825 ;
        RECT 51.055 35.655 51.345 35.825 ;
        RECT 51.515 35.655 51.805 35.825 ;
        RECT 51.975 35.655 52.265 35.825 ;
        RECT 52.435 35.655 52.725 35.825 ;
        RECT 52.895 35.655 53.185 35.825 ;
        RECT 53.355 35.655 53.645 35.825 ;
        RECT 53.815 35.655 54.105 35.825 ;
        RECT 54.275 35.655 54.565 35.825 ;
        RECT 54.735 35.655 55.025 35.825 ;
        RECT 55.195 35.655 55.485 35.825 ;
        RECT 55.655 35.655 55.945 35.825 ;
        RECT 56.115 35.655 56.405 35.825 ;
        RECT 56.575 35.655 56.865 35.825 ;
        RECT 57.035 35.655 57.325 35.825 ;
        RECT 57.495 35.655 57.785 35.825 ;
        RECT 57.955 35.655 58.245 35.825 ;
        RECT 58.415 35.655 58.705 35.825 ;
        RECT 58.875 35.655 59.165 35.825 ;
        RECT 59.335 35.655 59.625 35.825 ;
        RECT 59.795 35.655 60.085 35.825 ;
        RECT 60.255 35.655 60.545 35.825 ;
        RECT 60.715 35.655 61.005 35.825 ;
        RECT 61.175 35.655 61.465 35.825 ;
        RECT 61.635 35.655 61.925 35.825 ;
        RECT 62.095 35.655 62.385 35.825 ;
        RECT 62.555 35.655 62.845 35.825 ;
        RECT 63.015 35.655 63.305 35.825 ;
        RECT 63.475 35.655 63.765 35.825 ;
        RECT 63.935 35.655 64.225 35.825 ;
        RECT 64.395 35.655 64.685 35.825 ;
        RECT 64.855 35.655 65.145 35.825 ;
        RECT 65.315 35.655 65.605 35.825 ;
        RECT 65.775 35.655 66.065 35.825 ;
        RECT 66.235 35.655 66.525 35.825 ;
        RECT 66.695 35.655 66.985 35.825 ;
        RECT 67.155 35.655 67.445 35.825 ;
        RECT 67.615 35.655 67.905 35.825 ;
        RECT 68.075 35.655 68.365 35.825 ;
        RECT 68.535 35.655 68.825 35.825 ;
        RECT 68.995 35.655 69.285 35.825 ;
        RECT 69.455 35.655 69.745 35.825 ;
        RECT 69.915 35.655 70.205 35.825 ;
        RECT 70.375 35.655 70.665 35.825 ;
        RECT 70.835 35.655 71.125 35.825 ;
        RECT 71.295 35.655 71.585 35.825 ;
        RECT 71.755 35.655 72.045 35.825 ;
        RECT 72.215 35.655 72.505 35.825 ;
        RECT 72.675 35.655 72.965 35.825 ;
        RECT 73.135 35.655 73.425 35.825 ;
        RECT 73.595 35.655 73.885 35.825 ;
        RECT 74.055 35.655 74.345 35.825 ;
        RECT 74.515 35.655 74.805 35.825 ;
        RECT 74.975 35.655 75.265 35.825 ;
        RECT 75.435 35.655 75.725 35.825 ;
        RECT 75.895 35.655 76.185 35.825 ;
        RECT 76.355 35.655 76.645 35.825 ;
        RECT 76.815 35.655 77.105 35.825 ;
        RECT 77.275 35.655 77.565 35.825 ;
        RECT 77.735 35.655 78.025 35.825 ;
        RECT 78.195 35.655 78.485 35.825 ;
        RECT 78.655 35.655 78.945 35.825 ;
        RECT 79.115 35.655 79.405 35.825 ;
        RECT 79.575 35.655 79.865 35.825 ;
        RECT 80.035 35.655 80.325 35.825 ;
        RECT 80.495 35.655 80.785 35.825 ;
        RECT 80.955 35.655 81.245 35.825 ;
        RECT 81.415 35.655 81.705 35.825 ;
        RECT 81.875 35.655 82.165 35.825 ;
        RECT 82.335 35.655 82.625 35.825 ;
        RECT 82.795 35.655 83.085 35.825 ;
        RECT 83.255 35.655 83.545 35.825 ;
        RECT 83.715 35.655 84.005 35.825 ;
        RECT 84.175 35.655 84.465 35.825 ;
        RECT 84.635 35.655 84.925 35.825 ;
        RECT 85.095 35.655 85.385 35.825 ;
        RECT 85.555 35.655 85.845 35.825 ;
        RECT 86.015 35.655 86.305 35.825 ;
        RECT 86.475 35.655 86.765 35.825 ;
        RECT 86.935 35.655 87.225 35.825 ;
        RECT 87.395 35.655 87.685 35.825 ;
        RECT 87.855 35.655 88.145 35.825 ;
        RECT 88.315 35.655 88.605 35.825 ;
        RECT 88.775 35.655 89.065 35.825 ;
        RECT 89.235 35.655 89.525 35.825 ;
        RECT 89.695 35.655 89.985 35.825 ;
        RECT 90.155 35.655 90.445 35.825 ;
        RECT 90.615 35.655 90.905 35.825 ;
        RECT 91.075 35.655 91.365 35.825 ;
        RECT 91.535 35.655 91.825 35.825 ;
        RECT 91.995 35.655 92.285 35.825 ;
        RECT 92.455 35.655 92.745 35.825 ;
        RECT 92.915 35.655 93.205 35.825 ;
        RECT 93.375 35.655 93.665 35.825 ;
        RECT 93.835 35.655 94.125 35.825 ;
        RECT 94.295 35.655 94.585 35.825 ;
        RECT 94.755 35.655 95.045 35.825 ;
        RECT 95.215 35.655 95.505 35.825 ;
        RECT 95.675 35.655 95.965 35.825 ;
        RECT 96.135 35.655 96.425 35.825 ;
        RECT 96.595 35.655 96.885 35.825 ;
        RECT 97.055 35.655 97.345 35.825 ;
        RECT 97.515 35.655 97.805 35.825 ;
        RECT 97.975 35.655 98.265 35.825 ;
        RECT 98.435 35.655 98.725 35.825 ;
        RECT 98.895 35.655 99.185 35.825 ;
        RECT 99.355 35.655 99.645 35.825 ;
        RECT 99.815 35.655 99.960 35.825 ;
        RECT 16.785 34.905 17.995 35.655 ;
        RECT 18.165 34.905 19.375 35.655 ;
        RECT 16.785 34.365 17.305 34.905 ;
        RECT 17.475 34.195 17.995 34.735 ;
        RECT 18.165 34.365 18.685 34.905 ;
        RECT 18.855 34.195 19.375 34.735 ;
        RECT 16.785 33.105 17.995 34.195 ;
        RECT 18.165 33.105 19.375 34.195 ;
      LAYER li1 ;
        RECT 19.545 34.000 20.065 35.485 ;
      LAYER li1 ;
        RECT 20.235 34.995 20.575 35.655 ;
        RECT 20.925 34.885 26.270 35.655 ;
        RECT 26.445 34.885 29.955 35.655 ;
        RECT 31.045 34.930 31.335 35.655 ;
        RECT 31.505 34.885 36.850 35.655 ;
        RECT 37.025 34.885 42.370 35.655 ;
        RECT 42.545 34.885 47.890 35.655 ;
        RECT 48.065 34.885 53.410 35.655 ;
        RECT 53.585 34.885 58.930 35.655 ;
        RECT 59.105 34.930 59.395 35.655 ;
        RECT 59.565 34.885 64.910 35.655 ;
        RECT 65.085 34.885 70.430 35.655 ;
        RECT 70.605 34.885 75.950 35.655 ;
        RECT 76.125 34.885 81.470 35.655 ;
        RECT 81.645 34.885 86.990 35.655 ;
        RECT 87.165 34.930 87.455 35.655 ;
        RECT 87.625 34.885 92.970 35.655 ;
        RECT 93.145 34.885 98.490 35.655 ;
        RECT 98.665 34.905 99.875 35.655 ;
        RECT 20.925 34.365 23.505 34.885 ;
        RECT 23.675 34.195 26.270 34.715 ;
        RECT 26.445 34.365 28.095 34.885 ;
        RECT 28.265 34.195 29.955 34.715 ;
        RECT 31.505 34.365 34.085 34.885 ;
        RECT 19.735 33.105 20.065 33.830 ;
        RECT 20.925 33.105 26.270 34.195 ;
        RECT 26.445 33.105 29.955 34.195 ;
        RECT 31.045 33.105 31.335 34.270 ;
        RECT 34.255 34.195 36.850 34.715 ;
        RECT 37.025 34.365 39.605 34.885 ;
        RECT 39.775 34.195 42.370 34.715 ;
        RECT 42.545 34.365 45.125 34.885 ;
        RECT 45.295 34.195 47.890 34.715 ;
        RECT 48.065 34.365 50.645 34.885 ;
        RECT 50.815 34.195 53.410 34.715 ;
        RECT 53.585 34.365 56.165 34.885 ;
        RECT 56.335 34.195 58.930 34.715 ;
        RECT 59.565 34.365 62.145 34.885 ;
        RECT 31.505 33.105 36.850 34.195 ;
        RECT 37.025 33.105 42.370 34.195 ;
        RECT 42.545 33.105 47.890 34.195 ;
        RECT 48.065 33.105 53.410 34.195 ;
        RECT 53.585 33.105 58.930 34.195 ;
        RECT 59.105 33.105 59.395 34.270 ;
        RECT 62.315 34.195 64.910 34.715 ;
        RECT 65.085 34.365 67.665 34.885 ;
        RECT 67.835 34.195 70.430 34.715 ;
        RECT 70.605 34.365 73.185 34.885 ;
        RECT 73.355 34.195 75.950 34.715 ;
        RECT 76.125 34.365 78.705 34.885 ;
        RECT 78.875 34.195 81.470 34.715 ;
        RECT 81.645 34.365 84.225 34.885 ;
        RECT 84.395 34.195 86.990 34.715 ;
        RECT 87.625 34.365 90.205 34.885 ;
        RECT 59.565 33.105 64.910 34.195 ;
        RECT 65.085 33.105 70.430 34.195 ;
        RECT 70.605 33.105 75.950 34.195 ;
        RECT 76.125 33.105 81.470 34.195 ;
        RECT 81.645 33.105 86.990 34.195 ;
        RECT 87.165 33.105 87.455 34.270 ;
        RECT 90.375 34.195 92.970 34.715 ;
        RECT 93.145 34.365 95.725 34.885 ;
        RECT 95.895 34.195 98.490 34.715 ;
        RECT 87.625 33.105 92.970 34.195 ;
        RECT 93.145 33.105 98.490 34.195 ;
        RECT 98.665 34.195 99.185 34.735 ;
        RECT 99.355 34.365 99.875 34.905 ;
        RECT 98.665 33.105 99.875 34.195 ;
        RECT 16.700 32.935 16.845 33.105 ;
        RECT 17.015 32.935 17.305 33.105 ;
        RECT 17.475 32.935 17.765 33.105 ;
        RECT 17.935 32.935 18.225 33.105 ;
        RECT 18.395 32.935 18.685 33.105 ;
        RECT 18.855 32.935 19.145 33.105 ;
        RECT 19.315 32.935 19.605 33.105 ;
        RECT 19.775 32.935 20.065 33.105 ;
        RECT 20.235 32.935 20.525 33.105 ;
        RECT 20.695 32.935 20.985 33.105 ;
        RECT 21.155 32.935 21.445 33.105 ;
        RECT 21.615 32.935 21.905 33.105 ;
        RECT 22.075 32.935 22.365 33.105 ;
        RECT 22.535 32.935 22.825 33.105 ;
        RECT 22.995 32.935 23.285 33.105 ;
        RECT 23.455 32.935 23.745 33.105 ;
        RECT 23.915 32.935 24.205 33.105 ;
        RECT 24.375 32.935 24.665 33.105 ;
        RECT 24.835 32.935 25.125 33.105 ;
        RECT 25.295 32.935 25.585 33.105 ;
        RECT 25.755 32.935 26.045 33.105 ;
        RECT 26.215 32.935 26.505 33.105 ;
        RECT 26.675 32.935 26.965 33.105 ;
        RECT 27.135 32.935 27.425 33.105 ;
        RECT 27.595 32.935 27.885 33.105 ;
        RECT 28.055 32.935 28.345 33.105 ;
        RECT 28.515 32.935 28.805 33.105 ;
        RECT 28.975 32.935 29.265 33.105 ;
        RECT 29.435 32.935 29.725 33.105 ;
        RECT 29.895 32.935 30.185 33.105 ;
        RECT 30.355 32.935 30.645 33.105 ;
        RECT 30.815 32.935 31.105 33.105 ;
        RECT 31.275 32.935 31.565 33.105 ;
        RECT 31.735 32.935 32.025 33.105 ;
        RECT 32.195 32.935 32.485 33.105 ;
        RECT 32.655 32.935 32.945 33.105 ;
        RECT 33.115 32.935 33.405 33.105 ;
        RECT 33.575 32.935 33.865 33.105 ;
        RECT 34.035 32.935 34.325 33.105 ;
        RECT 34.495 32.935 34.785 33.105 ;
        RECT 34.955 32.935 35.245 33.105 ;
        RECT 35.415 32.935 35.705 33.105 ;
        RECT 35.875 32.935 36.165 33.105 ;
        RECT 36.335 32.935 36.625 33.105 ;
        RECT 36.795 32.935 37.085 33.105 ;
        RECT 37.255 32.935 37.545 33.105 ;
        RECT 37.715 32.935 38.005 33.105 ;
        RECT 38.175 32.935 38.465 33.105 ;
        RECT 38.635 32.935 38.925 33.105 ;
        RECT 39.095 32.935 39.385 33.105 ;
        RECT 39.555 32.935 39.845 33.105 ;
        RECT 40.015 32.935 40.305 33.105 ;
        RECT 40.475 32.935 40.765 33.105 ;
        RECT 40.935 32.935 41.225 33.105 ;
        RECT 41.395 32.935 41.685 33.105 ;
        RECT 41.855 32.935 42.145 33.105 ;
        RECT 42.315 32.935 42.605 33.105 ;
        RECT 42.775 32.935 43.065 33.105 ;
        RECT 43.235 32.935 43.525 33.105 ;
        RECT 43.695 32.935 43.985 33.105 ;
        RECT 44.155 32.935 44.445 33.105 ;
        RECT 44.615 32.935 44.905 33.105 ;
        RECT 45.075 32.935 45.365 33.105 ;
        RECT 45.535 32.935 45.825 33.105 ;
        RECT 45.995 32.935 46.285 33.105 ;
        RECT 46.455 32.935 46.745 33.105 ;
        RECT 46.915 32.935 47.205 33.105 ;
        RECT 47.375 32.935 47.665 33.105 ;
        RECT 47.835 32.935 48.125 33.105 ;
        RECT 48.295 32.935 48.585 33.105 ;
        RECT 48.755 32.935 49.045 33.105 ;
        RECT 49.215 32.935 49.505 33.105 ;
        RECT 49.675 32.935 49.965 33.105 ;
        RECT 50.135 32.935 50.425 33.105 ;
        RECT 50.595 32.935 50.885 33.105 ;
        RECT 51.055 32.935 51.345 33.105 ;
        RECT 51.515 32.935 51.805 33.105 ;
        RECT 51.975 32.935 52.265 33.105 ;
        RECT 52.435 32.935 52.725 33.105 ;
        RECT 52.895 32.935 53.185 33.105 ;
        RECT 53.355 32.935 53.645 33.105 ;
        RECT 53.815 32.935 54.105 33.105 ;
        RECT 54.275 32.935 54.565 33.105 ;
        RECT 54.735 32.935 55.025 33.105 ;
        RECT 55.195 32.935 55.485 33.105 ;
        RECT 55.655 32.935 55.945 33.105 ;
        RECT 56.115 32.935 56.405 33.105 ;
        RECT 56.575 32.935 56.865 33.105 ;
        RECT 57.035 32.935 57.325 33.105 ;
        RECT 57.495 32.935 57.785 33.105 ;
        RECT 57.955 32.935 58.245 33.105 ;
        RECT 58.415 32.935 58.705 33.105 ;
        RECT 58.875 32.935 59.165 33.105 ;
        RECT 59.335 32.935 59.625 33.105 ;
        RECT 59.795 32.935 60.085 33.105 ;
        RECT 60.255 32.935 60.545 33.105 ;
        RECT 60.715 32.935 61.005 33.105 ;
        RECT 61.175 32.935 61.465 33.105 ;
        RECT 61.635 32.935 61.925 33.105 ;
        RECT 62.095 32.935 62.385 33.105 ;
        RECT 62.555 32.935 62.845 33.105 ;
        RECT 63.015 32.935 63.305 33.105 ;
        RECT 63.475 32.935 63.765 33.105 ;
        RECT 63.935 32.935 64.225 33.105 ;
        RECT 64.395 32.935 64.685 33.105 ;
        RECT 64.855 32.935 65.145 33.105 ;
        RECT 65.315 32.935 65.605 33.105 ;
        RECT 65.775 32.935 66.065 33.105 ;
        RECT 66.235 32.935 66.525 33.105 ;
        RECT 66.695 32.935 66.985 33.105 ;
        RECT 67.155 32.935 67.445 33.105 ;
        RECT 67.615 32.935 67.905 33.105 ;
        RECT 68.075 32.935 68.365 33.105 ;
        RECT 68.535 32.935 68.825 33.105 ;
        RECT 68.995 32.935 69.285 33.105 ;
        RECT 69.455 32.935 69.745 33.105 ;
        RECT 69.915 32.935 70.205 33.105 ;
        RECT 70.375 32.935 70.665 33.105 ;
        RECT 70.835 32.935 71.125 33.105 ;
        RECT 71.295 32.935 71.585 33.105 ;
        RECT 71.755 32.935 72.045 33.105 ;
        RECT 72.215 32.935 72.505 33.105 ;
        RECT 72.675 32.935 72.965 33.105 ;
        RECT 73.135 32.935 73.425 33.105 ;
        RECT 73.595 32.935 73.885 33.105 ;
        RECT 74.055 32.935 74.345 33.105 ;
        RECT 74.515 32.935 74.805 33.105 ;
        RECT 74.975 32.935 75.265 33.105 ;
        RECT 75.435 32.935 75.725 33.105 ;
        RECT 75.895 32.935 76.185 33.105 ;
        RECT 76.355 32.935 76.645 33.105 ;
        RECT 76.815 32.935 77.105 33.105 ;
        RECT 77.275 32.935 77.565 33.105 ;
        RECT 77.735 32.935 78.025 33.105 ;
        RECT 78.195 32.935 78.485 33.105 ;
        RECT 78.655 32.935 78.945 33.105 ;
        RECT 79.115 32.935 79.405 33.105 ;
        RECT 79.575 32.935 79.865 33.105 ;
        RECT 80.035 32.935 80.325 33.105 ;
        RECT 80.495 32.935 80.785 33.105 ;
        RECT 80.955 32.935 81.245 33.105 ;
        RECT 81.415 32.935 81.705 33.105 ;
        RECT 81.875 32.935 82.165 33.105 ;
        RECT 82.335 32.935 82.625 33.105 ;
        RECT 82.795 32.935 83.085 33.105 ;
        RECT 83.255 32.935 83.545 33.105 ;
        RECT 83.715 32.935 84.005 33.105 ;
        RECT 84.175 32.935 84.465 33.105 ;
        RECT 84.635 32.935 84.925 33.105 ;
        RECT 85.095 32.935 85.385 33.105 ;
        RECT 85.555 32.935 85.845 33.105 ;
        RECT 86.015 32.935 86.305 33.105 ;
        RECT 86.475 32.935 86.765 33.105 ;
        RECT 86.935 32.935 87.225 33.105 ;
        RECT 87.395 32.935 87.685 33.105 ;
        RECT 87.855 32.935 88.145 33.105 ;
        RECT 88.315 32.935 88.605 33.105 ;
        RECT 88.775 32.935 89.065 33.105 ;
        RECT 89.235 32.935 89.525 33.105 ;
        RECT 89.695 32.935 89.985 33.105 ;
        RECT 90.155 32.935 90.445 33.105 ;
        RECT 90.615 32.935 90.905 33.105 ;
        RECT 91.075 32.935 91.365 33.105 ;
        RECT 91.535 32.935 91.825 33.105 ;
        RECT 91.995 32.935 92.285 33.105 ;
        RECT 92.455 32.935 92.745 33.105 ;
        RECT 92.915 32.935 93.205 33.105 ;
        RECT 93.375 32.935 93.665 33.105 ;
        RECT 93.835 32.935 94.125 33.105 ;
        RECT 94.295 32.935 94.585 33.105 ;
        RECT 94.755 32.935 95.045 33.105 ;
        RECT 95.215 32.935 95.505 33.105 ;
        RECT 95.675 32.935 95.965 33.105 ;
        RECT 96.135 32.935 96.425 33.105 ;
        RECT 96.595 32.935 96.885 33.105 ;
        RECT 97.055 32.935 97.345 33.105 ;
        RECT 97.515 32.935 97.805 33.105 ;
        RECT 97.975 32.935 98.265 33.105 ;
        RECT 98.435 32.935 98.725 33.105 ;
        RECT 98.895 32.935 99.185 33.105 ;
        RECT 99.355 32.935 99.645 33.105 ;
        RECT 99.815 32.935 99.960 33.105 ;
        RECT 16.785 31.845 17.995 32.935 ;
        RECT 18.165 31.845 23.510 32.935 ;
        RECT 23.685 31.845 29.030 32.935 ;
        RECT 29.205 31.845 34.550 32.935 ;
        RECT 34.725 31.845 40.070 32.935 ;
        RECT 40.245 31.845 43.755 32.935 ;
        RECT 16.785 31.135 17.305 31.675 ;
        RECT 17.475 31.305 17.995 31.845 ;
        RECT 18.165 31.155 20.745 31.675 ;
        RECT 20.915 31.325 23.510 31.845 ;
        RECT 23.685 31.155 26.265 31.675 ;
        RECT 26.435 31.325 29.030 31.845 ;
        RECT 29.205 31.155 31.785 31.675 ;
        RECT 31.955 31.325 34.550 31.845 ;
        RECT 34.725 31.155 37.305 31.675 ;
        RECT 37.475 31.325 40.070 31.845 ;
        RECT 40.245 31.155 41.895 31.675 ;
        RECT 42.065 31.325 43.755 31.845 ;
        RECT 44.845 31.770 45.135 32.935 ;
        RECT 45.305 31.845 50.650 32.935 ;
        RECT 50.825 31.845 56.170 32.935 ;
        RECT 56.345 31.845 61.690 32.935 ;
        RECT 61.865 31.845 67.210 32.935 ;
        RECT 67.385 31.845 72.730 32.935 ;
        RECT 45.305 31.155 47.885 31.675 ;
        RECT 48.055 31.325 50.650 31.845 ;
        RECT 50.825 31.155 53.405 31.675 ;
        RECT 53.575 31.325 56.170 31.845 ;
        RECT 56.345 31.155 58.925 31.675 ;
        RECT 59.095 31.325 61.690 31.845 ;
        RECT 61.865 31.155 64.445 31.675 ;
        RECT 64.615 31.325 67.210 31.845 ;
        RECT 67.385 31.155 69.965 31.675 ;
        RECT 70.135 31.325 72.730 31.845 ;
        RECT 72.905 31.770 73.195 32.935 ;
        RECT 73.365 31.845 78.710 32.935 ;
        RECT 78.885 31.845 84.230 32.935 ;
        RECT 84.405 31.845 89.750 32.935 ;
        RECT 89.925 31.845 95.270 32.935 ;
        RECT 95.445 31.845 98.035 32.935 ;
        RECT 73.365 31.155 75.945 31.675 ;
        RECT 76.115 31.325 78.710 31.845 ;
        RECT 78.885 31.155 81.465 31.675 ;
        RECT 81.635 31.325 84.230 31.845 ;
        RECT 84.405 31.155 86.985 31.675 ;
        RECT 87.155 31.325 89.750 31.845 ;
        RECT 89.925 31.155 92.505 31.675 ;
        RECT 92.675 31.325 95.270 31.845 ;
        RECT 95.445 31.155 96.655 31.675 ;
        RECT 96.825 31.325 98.035 31.845 ;
        RECT 98.665 31.845 99.875 32.935 ;
        RECT 98.665 31.305 99.185 31.845 ;
        RECT 16.785 30.385 17.995 31.135 ;
        RECT 18.165 30.385 23.510 31.155 ;
        RECT 23.685 30.385 29.030 31.155 ;
        RECT 29.205 30.385 34.550 31.155 ;
        RECT 34.725 30.385 40.070 31.155 ;
        RECT 40.245 30.385 43.755 31.155 ;
        RECT 44.845 30.385 45.135 31.110 ;
        RECT 45.305 30.385 50.650 31.155 ;
        RECT 50.825 30.385 56.170 31.155 ;
        RECT 56.345 30.385 61.690 31.155 ;
        RECT 61.865 30.385 67.210 31.155 ;
        RECT 67.385 30.385 72.730 31.155 ;
        RECT 72.905 30.385 73.195 31.110 ;
        RECT 73.365 30.385 78.710 31.155 ;
        RECT 78.885 30.385 84.230 31.155 ;
        RECT 84.405 30.385 89.750 31.155 ;
        RECT 89.925 30.385 95.270 31.155 ;
        RECT 95.445 30.385 98.035 31.155 ;
        RECT 99.355 31.135 99.875 31.675 ;
        RECT 98.665 30.385 99.875 31.135 ;
        RECT 16.700 30.215 16.845 30.385 ;
        RECT 17.015 30.215 17.305 30.385 ;
        RECT 17.475 30.215 17.765 30.385 ;
        RECT 17.935 30.215 18.225 30.385 ;
        RECT 18.395 30.215 18.685 30.385 ;
        RECT 18.855 30.215 19.145 30.385 ;
        RECT 19.315 30.215 19.605 30.385 ;
        RECT 19.775 30.215 20.065 30.385 ;
        RECT 20.235 30.215 20.525 30.385 ;
        RECT 20.695 30.215 20.985 30.385 ;
        RECT 21.155 30.215 21.445 30.385 ;
        RECT 21.615 30.215 21.905 30.385 ;
        RECT 22.075 30.215 22.365 30.385 ;
        RECT 22.535 30.215 22.825 30.385 ;
        RECT 22.995 30.215 23.285 30.385 ;
        RECT 23.455 30.215 23.745 30.385 ;
        RECT 23.915 30.215 24.205 30.385 ;
        RECT 24.375 30.215 24.665 30.385 ;
        RECT 24.835 30.215 25.125 30.385 ;
        RECT 25.295 30.215 25.585 30.385 ;
        RECT 25.755 30.215 26.045 30.385 ;
        RECT 26.215 30.215 26.505 30.385 ;
        RECT 26.675 30.215 26.965 30.385 ;
        RECT 27.135 30.215 27.425 30.385 ;
        RECT 27.595 30.215 27.885 30.385 ;
        RECT 28.055 30.215 28.345 30.385 ;
        RECT 28.515 30.215 28.805 30.385 ;
        RECT 28.975 30.215 29.265 30.385 ;
        RECT 29.435 30.215 29.725 30.385 ;
        RECT 29.895 30.215 30.185 30.385 ;
        RECT 30.355 30.215 30.645 30.385 ;
        RECT 30.815 30.215 31.105 30.385 ;
        RECT 31.275 30.215 31.565 30.385 ;
        RECT 31.735 30.215 32.025 30.385 ;
        RECT 32.195 30.215 32.485 30.385 ;
        RECT 32.655 30.215 32.945 30.385 ;
        RECT 33.115 30.215 33.405 30.385 ;
        RECT 33.575 30.215 33.865 30.385 ;
        RECT 34.035 30.215 34.325 30.385 ;
        RECT 34.495 30.215 34.785 30.385 ;
        RECT 34.955 30.215 35.245 30.385 ;
        RECT 35.415 30.215 35.705 30.385 ;
        RECT 35.875 30.215 36.165 30.385 ;
        RECT 36.335 30.215 36.625 30.385 ;
        RECT 36.795 30.215 37.085 30.385 ;
        RECT 37.255 30.215 37.545 30.385 ;
        RECT 37.715 30.215 38.005 30.385 ;
        RECT 38.175 30.215 38.465 30.385 ;
        RECT 38.635 30.215 38.925 30.385 ;
        RECT 39.095 30.215 39.385 30.385 ;
        RECT 39.555 30.215 39.845 30.385 ;
        RECT 40.015 30.215 40.305 30.385 ;
        RECT 40.475 30.215 40.765 30.385 ;
        RECT 40.935 30.215 41.225 30.385 ;
        RECT 41.395 30.215 41.685 30.385 ;
        RECT 41.855 30.215 42.145 30.385 ;
        RECT 42.315 30.215 42.605 30.385 ;
        RECT 42.775 30.215 43.065 30.385 ;
        RECT 43.235 30.215 43.525 30.385 ;
        RECT 43.695 30.215 43.985 30.385 ;
        RECT 44.155 30.215 44.445 30.385 ;
        RECT 44.615 30.215 44.905 30.385 ;
        RECT 45.075 30.215 45.365 30.385 ;
        RECT 45.535 30.215 45.825 30.385 ;
        RECT 45.995 30.215 46.285 30.385 ;
        RECT 46.455 30.215 46.745 30.385 ;
        RECT 46.915 30.215 47.205 30.385 ;
        RECT 47.375 30.215 47.665 30.385 ;
        RECT 47.835 30.215 48.125 30.385 ;
        RECT 48.295 30.215 48.585 30.385 ;
        RECT 48.755 30.215 49.045 30.385 ;
        RECT 49.215 30.215 49.505 30.385 ;
        RECT 49.675 30.215 49.965 30.385 ;
        RECT 50.135 30.215 50.425 30.385 ;
        RECT 50.595 30.215 50.885 30.385 ;
        RECT 51.055 30.215 51.345 30.385 ;
        RECT 51.515 30.215 51.805 30.385 ;
        RECT 51.975 30.215 52.265 30.385 ;
        RECT 52.435 30.215 52.725 30.385 ;
        RECT 52.895 30.215 53.185 30.385 ;
        RECT 53.355 30.215 53.645 30.385 ;
        RECT 53.815 30.215 54.105 30.385 ;
        RECT 54.275 30.215 54.565 30.385 ;
        RECT 54.735 30.215 55.025 30.385 ;
        RECT 55.195 30.215 55.485 30.385 ;
        RECT 55.655 30.215 55.945 30.385 ;
        RECT 56.115 30.215 56.405 30.385 ;
        RECT 56.575 30.215 56.865 30.385 ;
        RECT 57.035 30.215 57.325 30.385 ;
        RECT 57.495 30.215 57.785 30.385 ;
        RECT 57.955 30.215 58.245 30.385 ;
        RECT 58.415 30.215 58.705 30.385 ;
        RECT 58.875 30.215 59.165 30.385 ;
        RECT 59.335 30.215 59.625 30.385 ;
        RECT 59.795 30.215 60.085 30.385 ;
        RECT 60.255 30.215 60.545 30.385 ;
        RECT 60.715 30.215 61.005 30.385 ;
        RECT 61.175 30.215 61.465 30.385 ;
        RECT 61.635 30.215 61.925 30.385 ;
        RECT 62.095 30.215 62.385 30.385 ;
        RECT 62.555 30.215 62.845 30.385 ;
        RECT 63.015 30.215 63.305 30.385 ;
        RECT 63.475 30.215 63.765 30.385 ;
        RECT 63.935 30.215 64.225 30.385 ;
        RECT 64.395 30.215 64.685 30.385 ;
        RECT 64.855 30.215 65.145 30.385 ;
        RECT 65.315 30.215 65.605 30.385 ;
        RECT 65.775 30.215 66.065 30.385 ;
        RECT 66.235 30.215 66.525 30.385 ;
        RECT 66.695 30.215 66.985 30.385 ;
        RECT 67.155 30.215 67.445 30.385 ;
        RECT 67.615 30.215 67.905 30.385 ;
        RECT 68.075 30.215 68.365 30.385 ;
        RECT 68.535 30.215 68.825 30.385 ;
        RECT 68.995 30.215 69.285 30.385 ;
        RECT 69.455 30.215 69.745 30.385 ;
        RECT 69.915 30.215 70.205 30.385 ;
        RECT 70.375 30.215 70.665 30.385 ;
        RECT 70.835 30.215 71.125 30.385 ;
        RECT 71.295 30.215 71.585 30.385 ;
        RECT 71.755 30.215 72.045 30.385 ;
        RECT 72.215 30.215 72.505 30.385 ;
        RECT 72.675 30.215 72.965 30.385 ;
        RECT 73.135 30.215 73.425 30.385 ;
        RECT 73.595 30.215 73.885 30.385 ;
        RECT 74.055 30.215 74.345 30.385 ;
        RECT 74.515 30.215 74.805 30.385 ;
        RECT 74.975 30.215 75.265 30.385 ;
        RECT 75.435 30.215 75.725 30.385 ;
        RECT 75.895 30.215 76.185 30.385 ;
        RECT 76.355 30.215 76.645 30.385 ;
        RECT 76.815 30.215 77.105 30.385 ;
        RECT 77.275 30.215 77.565 30.385 ;
        RECT 77.735 30.215 78.025 30.385 ;
        RECT 78.195 30.215 78.485 30.385 ;
        RECT 78.655 30.215 78.945 30.385 ;
        RECT 79.115 30.215 79.405 30.385 ;
        RECT 79.575 30.215 79.865 30.385 ;
        RECT 80.035 30.215 80.325 30.385 ;
        RECT 80.495 30.215 80.785 30.385 ;
        RECT 80.955 30.215 81.245 30.385 ;
        RECT 81.415 30.215 81.705 30.385 ;
        RECT 81.875 30.215 82.165 30.385 ;
        RECT 82.335 30.215 82.625 30.385 ;
        RECT 82.795 30.215 83.085 30.385 ;
        RECT 83.255 30.215 83.545 30.385 ;
        RECT 83.715 30.215 84.005 30.385 ;
        RECT 84.175 30.215 84.465 30.385 ;
        RECT 84.635 30.215 84.925 30.385 ;
        RECT 85.095 30.215 85.385 30.385 ;
        RECT 85.555 30.215 85.845 30.385 ;
        RECT 86.015 30.215 86.305 30.385 ;
        RECT 86.475 30.215 86.765 30.385 ;
        RECT 86.935 30.215 87.225 30.385 ;
        RECT 87.395 30.215 87.685 30.385 ;
        RECT 87.855 30.215 88.145 30.385 ;
        RECT 88.315 30.215 88.605 30.385 ;
        RECT 88.775 30.215 89.065 30.385 ;
        RECT 89.235 30.215 89.525 30.385 ;
        RECT 89.695 30.215 89.985 30.385 ;
        RECT 90.155 30.215 90.445 30.385 ;
        RECT 90.615 30.215 90.905 30.385 ;
        RECT 91.075 30.215 91.365 30.385 ;
        RECT 91.535 30.215 91.825 30.385 ;
        RECT 91.995 30.215 92.285 30.385 ;
        RECT 92.455 30.215 92.745 30.385 ;
        RECT 92.915 30.215 93.205 30.385 ;
        RECT 93.375 30.215 93.665 30.385 ;
        RECT 93.835 30.215 94.125 30.385 ;
        RECT 94.295 30.215 94.585 30.385 ;
        RECT 94.755 30.215 95.045 30.385 ;
        RECT 95.215 30.215 95.505 30.385 ;
        RECT 95.675 30.215 95.965 30.385 ;
        RECT 96.135 30.215 96.425 30.385 ;
        RECT 96.595 30.215 96.885 30.385 ;
        RECT 97.055 30.215 97.345 30.385 ;
        RECT 97.515 30.215 97.805 30.385 ;
        RECT 97.975 30.215 98.265 30.385 ;
        RECT 98.435 30.215 98.725 30.385 ;
        RECT 98.895 30.215 99.185 30.385 ;
        RECT 99.355 30.215 99.645 30.385 ;
        RECT 99.815 30.215 99.960 30.385 ;
        RECT 16.785 29.465 17.995 30.215 ;
        RECT 16.785 28.925 17.305 29.465 ;
        RECT 18.165 29.445 23.510 30.215 ;
        RECT 23.685 29.445 29.030 30.215 ;
        RECT 29.205 29.445 30.875 30.215 ;
        RECT 31.045 29.490 31.335 30.215 ;
        RECT 31.505 29.445 36.850 30.215 ;
        RECT 37.025 29.445 42.370 30.215 ;
        RECT 42.545 29.445 47.890 30.215 ;
        RECT 48.065 29.445 53.410 30.215 ;
        RECT 53.585 29.445 58.930 30.215 ;
        RECT 59.105 29.490 59.395 30.215 ;
        RECT 59.565 29.445 64.910 30.215 ;
        RECT 65.085 29.445 70.430 30.215 ;
        RECT 70.605 29.445 75.950 30.215 ;
        RECT 76.125 29.445 81.470 30.215 ;
        RECT 81.645 29.445 86.990 30.215 ;
        RECT 87.165 29.490 87.455 30.215 ;
        RECT 87.625 29.445 92.970 30.215 ;
        RECT 93.145 29.445 98.490 30.215 ;
        RECT 98.665 29.465 99.875 30.215 ;
        RECT 17.475 28.755 17.995 29.295 ;
        RECT 18.165 28.925 20.745 29.445 ;
        RECT 20.915 28.755 23.510 29.275 ;
        RECT 23.685 28.925 26.265 29.445 ;
        RECT 26.435 28.755 29.030 29.275 ;
        RECT 29.205 28.925 29.955 29.445 ;
        RECT 30.125 28.755 30.875 29.275 ;
        RECT 31.505 28.925 34.085 29.445 ;
        RECT 16.785 27.665 17.995 28.755 ;
        RECT 18.165 27.665 23.510 28.755 ;
        RECT 23.685 27.665 29.030 28.755 ;
        RECT 29.205 27.665 30.875 28.755 ;
        RECT 31.045 27.665 31.335 28.830 ;
        RECT 34.255 28.755 36.850 29.275 ;
        RECT 37.025 28.925 39.605 29.445 ;
        RECT 39.775 28.755 42.370 29.275 ;
        RECT 42.545 28.925 45.125 29.445 ;
        RECT 45.295 28.755 47.890 29.275 ;
        RECT 48.065 28.925 50.645 29.445 ;
        RECT 50.815 28.755 53.410 29.275 ;
        RECT 53.585 28.925 56.165 29.445 ;
        RECT 56.335 28.755 58.930 29.275 ;
        RECT 59.565 28.925 62.145 29.445 ;
        RECT 31.505 27.665 36.850 28.755 ;
        RECT 37.025 27.665 42.370 28.755 ;
        RECT 42.545 27.665 47.890 28.755 ;
        RECT 48.065 27.665 53.410 28.755 ;
        RECT 53.585 27.665 58.930 28.755 ;
        RECT 59.105 27.665 59.395 28.830 ;
        RECT 62.315 28.755 64.910 29.275 ;
        RECT 65.085 28.925 67.665 29.445 ;
        RECT 67.835 28.755 70.430 29.275 ;
        RECT 70.605 28.925 73.185 29.445 ;
        RECT 73.355 28.755 75.950 29.275 ;
        RECT 76.125 28.925 78.705 29.445 ;
        RECT 78.875 28.755 81.470 29.275 ;
        RECT 81.645 28.925 84.225 29.445 ;
        RECT 84.395 28.755 86.990 29.275 ;
        RECT 87.625 28.925 90.205 29.445 ;
        RECT 59.565 27.665 64.910 28.755 ;
        RECT 65.085 27.665 70.430 28.755 ;
        RECT 70.605 27.665 75.950 28.755 ;
        RECT 76.125 27.665 81.470 28.755 ;
        RECT 81.645 27.665 86.990 28.755 ;
        RECT 87.165 27.665 87.455 28.830 ;
        RECT 90.375 28.755 92.970 29.275 ;
        RECT 93.145 28.925 95.725 29.445 ;
        RECT 95.895 28.755 98.490 29.275 ;
        RECT 87.625 27.665 92.970 28.755 ;
        RECT 93.145 27.665 98.490 28.755 ;
        RECT 98.665 28.755 99.185 29.295 ;
        RECT 99.355 28.925 99.875 29.465 ;
        RECT 98.665 27.665 99.875 28.755 ;
        RECT 16.700 27.495 16.845 27.665 ;
        RECT 17.015 27.495 17.305 27.665 ;
        RECT 17.475 27.495 17.765 27.665 ;
        RECT 17.935 27.495 18.225 27.665 ;
        RECT 18.395 27.495 18.685 27.665 ;
        RECT 18.855 27.495 19.145 27.665 ;
        RECT 19.315 27.495 19.605 27.665 ;
        RECT 19.775 27.495 20.065 27.665 ;
        RECT 20.235 27.495 20.525 27.665 ;
        RECT 20.695 27.495 20.985 27.665 ;
        RECT 21.155 27.495 21.445 27.665 ;
        RECT 21.615 27.495 21.905 27.665 ;
        RECT 22.075 27.495 22.365 27.665 ;
        RECT 22.535 27.495 22.825 27.665 ;
        RECT 22.995 27.495 23.285 27.665 ;
        RECT 23.455 27.495 23.745 27.665 ;
        RECT 23.915 27.495 24.205 27.665 ;
        RECT 24.375 27.495 24.665 27.665 ;
        RECT 24.835 27.495 25.125 27.665 ;
        RECT 25.295 27.495 25.585 27.665 ;
        RECT 25.755 27.495 26.045 27.665 ;
        RECT 26.215 27.495 26.505 27.665 ;
        RECT 26.675 27.495 26.965 27.665 ;
        RECT 27.135 27.495 27.425 27.665 ;
        RECT 27.595 27.495 27.885 27.665 ;
        RECT 28.055 27.495 28.345 27.665 ;
        RECT 28.515 27.495 28.805 27.665 ;
        RECT 28.975 27.495 29.265 27.665 ;
        RECT 29.435 27.495 29.725 27.665 ;
        RECT 29.895 27.495 30.185 27.665 ;
        RECT 30.355 27.495 30.645 27.665 ;
        RECT 30.815 27.495 31.105 27.665 ;
        RECT 31.275 27.495 31.565 27.665 ;
        RECT 31.735 27.495 32.025 27.665 ;
        RECT 32.195 27.495 32.485 27.665 ;
        RECT 32.655 27.495 32.945 27.665 ;
        RECT 33.115 27.495 33.405 27.665 ;
        RECT 33.575 27.495 33.865 27.665 ;
        RECT 34.035 27.495 34.325 27.665 ;
        RECT 34.495 27.495 34.785 27.665 ;
        RECT 34.955 27.495 35.245 27.665 ;
        RECT 35.415 27.495 35.705 27.665 ;
        RECT 35.875 27.495 36.165 27.665 ;
        RECT 36.335 27.495 36.625 27.665 ;
        RECT 36.795 27.495 37.085 27.665 ;
        RECT 37.255 27.495 37.545 27.665 ;
        RECT 37.715 27.495 38.005 27.665 ;
        RECT 38.175 27.495 38.465 27.665 ;
        RECT 38.635 27.495 38.925 27.665 ;
        RECT 39.095 27.495 39.385 27.665 ;
        RECT 39.555 27.495 39.845 27.665 ;
        RECT 40.015 27.495 40.305 27.665 ;
        RECT 40.475 27.495 40.765 27.665 ;
        RECT 40.935 27.495 41.225 27.665 ;
        RECT 41.395 27.495 41.685 27.665 ;
        RECT 41.855 27.495 42.145 27.665 ;
        RECT 42.315 27.495 42.605 27.665 ;
        RECT 42.775 27.495 43.065 27.665 ;
        RECT 43.235 27.495 43.525 27.665 ;
        RECT 43.695 27.495 43.985 27.665 ;
        RECT 44.155 27.495 44.445 27.665 ;
        RECT 44.615 27.495 44.905 27.665 ;
        RECT 45.075 27.495 45.365 27.665 ;
        RECT 45.535 27.495 45.825 27.665 ;
        RECT 45.995 27.495 46.285 27.665 ;
        RECT 46.455 27.495 46.745 27.665 ;
        RECT 46.915 27.495 47.205 27.665 ;
        RECT 47.375 27.495 47.665 27.665 ;
        RECT 47.835 27.495 48.125 27.665 ;
        RECT 48.295 27.495 48.585 27.665 ;
        RECT 48.755 27.495 49.045 27.665 ;
        RECT 49.215 27.495 49.505 27.665 ;
        RECT 49.675 27.495 49.965 27.665 ;
        RECT 50.135 27.495 50.425 27.665 ;
        RECT 50.595 27.495 50.885 27.665 ;
        RECT 51.055 27.495 51.345 27.665 ;
        RECT 51.515 27.495 51.805 27.665 ;
        RECT 51.975 27.495 52.265 27.665 ;
        RECT 52.435 27.495 52.725 27.665 ;
        RECT 52.895 27.495 53.185 27.665 ;
        RECT 53.355 27.495 53.645 27.665 ;
        RECT 53.815 27.495 54.105 27.665 ;
        RECT 54.275 27.495 54.565 27.665 ;
        RECT 54.735 27.495 55.025 27.665 ;
        RECT 55.195 27.495 55.485 27.665 ;
        RECT 55.655 27.495 55.945 27.665 ;
        RECT 56.115 27.495 56.405 27.665 ;
        RECT 56.575 27.495 56.865 27.665 ;
        RECT 57.035 27.495 57.325 27.665 ;
        RECT 57.495 27.495 57.785 27.665 ;
        RECT 57.955 27.495 58.245 27.665 ;
        RECT 58.415 27.495 58.705 27.665 ;
        RECT 58.875 27.495 59.165 27.665 ;
        RECT 59.335 27.495 59.625 27.665 ;
        RECT 59.795 27.495 60.085 27.665 ;
        RECT 60.255 27.495 60.545 27.665 ;
        RECT 60.715 27.495 61.005 27.665 ;
        RECT 61.175 27.495 61.465 27.665 ;
        RECT 61.635 27.495 61.925 27.665 ;
        RECT 62.095 27.495 62.385 27.665 ;
        RECT 62.555 27.495 62.845 27.665 ;
        RECT 63.015 27.495 63.305 27.665 ;
        RECT 63.475 27.495 63.765 27.665 ;
        RECT 63.935 27.495 64.225 27.665 ;
        RECT 64.395 27.495 64.685 27.665 ;
        RECT 64.855 27.495 65.145 27.665 ;
        RECT 65.315 27.495 65.605 27.665 ;
        RECT 65.775 27.495 66.065 27.665 ;
        RECT 66.235 27.495 66.525 27.665 ;
        RECT 66.695 27.495 66.985 27.665 ;
        RECT 67.155 27.495 67.445 27.665 ;
        RECT 67.615 27.495 67.905 27.665 ;
        RECT 68.075 27.495 68.365 27.665 ;
        RECT 68.535 27.495 68.825 27.665 ;
        RECT 68.995 27.495 69.285 27.665 ;
        RECT 69.455 27.495 69.745 27.665 ;
        RECT 69.915 27.495 70.205 27.665 ;
        RECT 70.375 27.495 70.665 27.665 ;
        RECT 70.835 27.495 71.125 27.665 ;
        RECT 71.295 27.495 71.585 27.665 ;
        RECT 71.755 27.495 72.045 27.665 ;
        RECT 72.215 27.495 72.505 27.665 ;
        RECT 72.675 27.495 72.965 27.665 ;
        RECT 73.135 27.495 73.425 27.665 ;
        RECT 73.595 27.495 73.885 27.665 ;
        RECT 74.055 27.495 74.345 27.665 ;
        RECT 74.515 27.495 74.805 27.665 ;
        RECT 74.975 27.495 75.265 27.665 ;
        RECT 75.435 27.495 75.725 27.665 ;
        RECT 75.895 27.495 76.185 27.665 ;
        RECT 76.355 27.495 76.645 27.665 ;
        RECT 76.815 27.495 77.105 27.665 ;
        RECT 77.275 27.495 77.565 27.665 ;
        RECT 77.735 27.495 78.025 27.665 ;
        RECT 78.195 27.495 78.485 27.665 ;
        RECT 78.655 27.495 78.945 27.665 ;
        RECT 79.115 27.495 79.405 27.665 ;
        RECT 79.575 27.495 79.865 27.665 ;
        RECT 80.035 27.495 80.325 27.665 ;
        RECT 80.495 27.495 80.785 27.665 ;
        RECT 80.955 27.495 81.245 27.665 ;
        RECT 81.415 27.495 81.705 27.665 ;
        RECT 81.875 27.495 82.165 27.665 ;
        RECT 82.335 27.495 82.625 27.665 ;
        RECT 82.795 27.495 83.085 27.665 ;
        RECT 83.255 27.495 83.545 27.665 ;
        RECT 83.715 27.495 84.005 27.665 ;
        RECT 84.175 27.495 84.465 27.665 ;
        RECT 84.635 27.495 84.925 27.665 ;
        RECT 85.095 27.495 85.385 27.665 ;
        RECT 85.555 27.495 85.845 27.665 ;
        RECT 86.015 27.495 86.305 27.665 ;
        RECT 86.475 27.495 86.765 27.665 ;
        RECT 86.935 27.495 87.225 27.665 ;
        RECT 87.395 27.495 87.685 27.665 ;
        RECT 87.855 27.495 88.145 27.665 ;
        RECT 88.315 27.495 88.605 27.665 ;
        RECT 88.775 27.495 89.065 27.665 ;
        RECT 89.235 27.495 89.525 27.665 ;
        RECT 89.695 27.495 89.985 27.665 ;
        RECT 90.155 27.495 90.445 27.665 ;
        RECT 90.615 27.495 90.905 27.665 ;
        RECT 91.075 27.495 91.365 27.665 ;
        RECT 91.535 27.495 91.825 27.665 ;
        RECT 91.995 27.495 92.285 27.665 ;
        RECT 92.455 27.495 92.745 27.665 ;
        RECT 92.915 27.495 93.205 27.665 ;
        RECT 93.375 27.495 93.665 27.665 ;
        RECT 93.835 27.495 94.125 27.665 ;
        RECT 94.295 27.495 94.585 27.665 ;
        RECT 94.755 27.495 95.045 27.665 ;
        RECT 95.215 27.495 95.505 27.665 ;
        RECT 95.675 27.495 95.965 27.665 ;
        RECT 96.135 27.495 96.425 27.665 ;
        RECT 96.595 27.495 96.885 27.665 ;
        RECT 97.055 27.495 97.345 27.665 ;
        RECT 97.515 27.495 97.805 27.665 ;
        RECT 97.975 27.495 98.265 27.665 ;
        RECT 98.435 27.495 98.725 27.665 ;
        RECT 98.895 27.495 99.185 27.665 ;
        RECT 99.355 27.495 99.645 27.665 ;
        RECT 99.815 27.495 99.960 27.665 ;
        RECT 16.785 26.405 17.995 27.495 ;
        RECT 18.165 26.405 23.510 27.495 ;
        RECT 23.685 26.405 29.030 27.495 ;
        RECT 29.205 26.405 34.550 27.495 ;
        RECT 34.725 26.405 40.070 27.495 ;
        RECT 40.245 26.405 43.755 27.495 ;
        RECT 16.785 25.695 17.305 26.235 ;
        RECT 17.475 25.865 17.995 26.405 ;
        RECT 18.165 25.715 20.745 26.235 ;
        RECT 20.915 25.885 23.510 26.405 ;
        RECT 23.685 25.715 26.265 26.235 ;
        RECT 26.435 25.885 29.030 26.405 ;
        RECT 29.205 25.715 31.785 26.235 ;
        RECT 31.955 25.885 34.550 26.405 ;
        RECT 34.725 25.715 37.305 26.235 ;
        RECT 37.475 25.885 40.070 26.405 ;
        RECT 40.245 25.715 41.895 26.235 ;
        RECT 42.065 25.885 43.755 26.405 ;
        RECT 44.845 26.330 45.135 27.495 ;
        RECT 45.305 26.405 50.650 27.495 ;
        RECT 50.825 26.405 56.170 27.495 ;
        RECT 56.345 26.405 61.690 27.495 ;
        RECT 61.865 26.405 67.210 27.495 ;
        RECT 67.385 26.405 72.730 27.495 ;
        RECT 45.305 25.715 47.885 26.235 ;
        RECT 48.055 25.885 50.650 26.405 ;
        RECT 50.825 25.715 53.405 26.235 ;
        RECT 53.575 25.885 56.170 26.405 ;
        RECT 56.345 25.715 58.925 26.235 ;
        RECT 59.095 25.885 61.690 26.405 ;
        RECT 61.865 25.715 64.445 26.235 ;
        RECT 64.615 25.885 67.210 26.405 ;
        RECT 67.385 25.715 69.965 26.235 ;
        RECT 70.135 25.885 72.730 26.405 ;
        RECT 72.905 26.330 73.195 27.495 ;
        RECT 73.365 26.405 78.710 27.495 ;
        RECT 78.885 26.405 84.230 27.495 ;
        RECT 84.405 26.405 89.750 27.495 ;
        RECT 89.925 26.405 95.270 27.495 ;
        RECT 95.445 26.405 98.035 27.495 ;
        RECT 73.365 25.715 75.945 26.235 ;
        RECT 76.115 25.885 78.710 26.405 ;
        RECT 78.885 25.715 81.465 26.235 ;
        RECT 81.635 25.885 84.230 26.405 ;
        RECT 84.405 25.715 86.985 26.235 ;
        RECT 87.155 25.885 89.750 26.405 ;
        RECT 89.925 25.715 92.505 26.235 ;
        RECT 92.675 25.885 95.270 26.405 ;
        RECT 95.445 25.715 96.655 26.235 ;
        RECT 96.825 25.885 98.035 26.405 ;
        RECT 98.665 26.405 99.875 27.495 ;
        RECT 98.665 25.865 99.185 26.405 ;
        RECT 16.785 24.945 17.995 25.695 ;
        RECT 18.165 24.945 23.510 25.715 ;
        RECT 23.685 24.945 29.030 25.715 ;
        RECT 29.205 24.945 34.550 25.715 ;
        RECT 34.725 24.945 40.070 25.715 ;
        RECT 40.245 24.945 43.755 25.715 ;
        RECT 44.845 24.945 45.135 25.670 ;
        RECT 45.305 24.945 50.650 25.715 ;
        RECT 50.825 24.945 56.170 25.715 ;
        RECT 56.345 24.945 61.690 25.715 ;
        RECT 61.865 24.945 67.210 25.715 ;
        RECT 67.385 24.945 72.730 25.715 ;
        RECT 72.905 24.945 73.195 25.670 ;
        RECT 73.365 24.945 78.710 25.715 ;
        RECT 78.885 24.945 84.230 25.715 ;
        RECT 84.405 24.945 89.750 25.715 ;
        RECT 89.925 24.945 95.270 25.715 ;
        RECT 95.445 24.945 98.035 25.715 ;
        RECT 99.355 25.695 99.875 26.235 ;
        RECT 98.665 24.945 99.875 25.695 ;
        RECT 16.700 24.775 16.845 24.945 ;
        RECT 17.015 24.775 17.305 24.945 ;
        RECT 17.475 24.775 17.765 24.945 ;
        RECT 17.935 24.775 18.225 24.945 ;
        RECT 18.395 24.775 18.685 24.945 ;
        RECT 18.855 24.775 19.145 24.945 ;
        RECT 19.315 24.775 19.605 24.945 ;
        RECT 19.775 24.775 20.065 24.945 ;
        RECT 20.235 24.775 20.525 24.945 ;
        RECT 20.695 24.775 20.985 24.945 ;
        RECT 21.155 24.775 21.445 24.945 ;
        RECT 21.615 24.775 21.905 24.945 ;
        RECT 22.075 24.775 22.365 24.945 ;
        RECT 22.535 24.775 22.825 24.945 ;
        RECT 22.995 24.775 23.285 24.945 ;
        RECT 23.455 24.775 23.745 24.945 ;
        RECT 23.915 24.775 24.205 24.945 ;
        RECT 24.375 24.775 24.665 24.945 ;
        RECT 24.835 24.775 25.125 24.945 ;
        RECT 25.295 24.775 25.585 24.945 ;
        RECT 25.755 24.775 26.045 24.945 ;
        RECT 26.215 24.775 26.505 24.945 ;
        RECT 26.675 24.775 26.965 24.945 ;
        RECT 27.135 24.775 27.425 24.945 ;
        RECT 27.595 24.775 27.885 24.945 ;
        RECT 28.055 24.775 28.345 24.945 ;
        RECT 28.515 24.775 28.805 24.945 ;
        RECT 28.975 24.775 29.265 24.945 ;
        RECT 29.435 24.775 29.725 24.945 ;
        RECT 29.895 24.775 30.185 24.945 ;
        RECT 30.355 24.775 30.645 24.945 ;
        RECT 30.815 24.775 31.105 24.945 ;
        RECT 31.275 24.775 31.565 24.945 ;
        RECT 31.735 24.775 32.025 24.945 ;
        RECT 32.195 24.775 32.485 24.945 ;
        RECT 32.655 24.775 32.945 24.945 ;
        RECT 33.115 24.775 33.405 24.945 ;
        RECT 33.575 24.775 33.865 24.945 ;
        RECT 34.035 24.775 34.325 24.945 ;
        RECT 34.495 24.775 34.785 24.945 ;
        RECT 34.955 24.775 35.245 24.945 ;
        RECT 35.415 24.775 35.705 24.945 ;
        RECT 35.875 24.775 36.165 24.945 ;
        RECT 36.335 24.775 36.625 24.945 ;
        RECT 36.795 24.775 37.085 24.945 ;
        RECT 37.255 24.775 37.545 24.945 ;
        RECT 37.715 24.775 38.005 24.945 ;
        RECT 38.175 24.775 38.465 24.945 ;
        RECT 38.635 24.775 38.925 24.945 ;
        RECT 39.095 24.775 39.385 24.945 ;
        RECT 39.555 24.775 39.845 24.945 ;
        RECT 40.015 24.775 40.305 24.945 ;
        RECT 40.475 24.775 40.765 24.945 ;
        RECT 40.935 24.775 41.225 24.945 ;
        RECT 41.395 24.775 41.685 24.945 ;
        RECT 41.855 24.775 42.145 24.945 ;
        RECT 42.315 24.775 42.605 24.945 ;
        RECT 42.775 24.775 43.065 24.945 ;
        RECT 43.235 24.775 43.525 24.945 ;
        RECT 43.695 24.775 43.985 24.945 ;
        RECT 44.155 24.775 44.445 24.945 ;
        RECT 44.615 24.775 44.905 24.945 ;
        RECT 45.075 24.775 45.365 24.945 ;
        RECT 45.535 24.775 45.825 24.945 ;
        RECT 45.995 24.775 46.285 24.945 ;
        RECT 46.455 24.775 46.745 24.945 ;
        RECT 46.915 24.775 47.205 24.945 ;
        RECT 47.375 24.775 47.665 24.945 ;
        RECT 47.835 24.775 48.125 24.945 ;
        RECT 48.295 24.775 48.585 24.945 ;
        RECT 48.755 24.775 49.045 24.945 ;
        RECT 49.215 24.775 49.505 24.945 ;
        RECT 49.675 24.775 49.965 24.945 ;
        RECT 50.135 24.775 50.425 24.945 ;
        RECT 50.595 24.775 50.885 24.945 ;
        RECT 51.055 24.775 51.345 24.945 ;
        RECT 51.515 24.775 51.805 24.945 ;
        RECT 51.975 24.775 52.265 24.945 ;
        RECT 52.435 24.775 52.725 24.945 ;
        RECT 52.895 24.775 53.185 24.945 ;
        RECT 53.355 24.775 53.645 24.945 ;
        RECT 53.815 24.775 54.105 24.945 ;
        RECT 54.275 24.775 54.565 24.945 ;
        RECT 54.735 24.775 55.025 24.945 ;
        RECT 55.195 24.775 55.485 24.945 ;
        RECT 55.655 24.775 55.945 24.945 ;
        RECT 56.115 24.775 56.405 24.945 ;
        RECT 56.575 24.775 56.865 24.945 ;
        RECT 57.035 24.775 57.325 24.945 ;
        RECT 57.495 24.775 57.785 24.945 ;
        RECT 57.955 24.775 58.245 24.945 ;
        RECT 58.415 24.775 58.705 24.945 ;
        RECT 58.875 24.775 59.165 24.945 ;
        RECT 59.335 24.775 59.625 24.945 ;
        RECT 59.795 24.775 60.085 24.945 ;
        RECT 60.255 24.775 60.545 24.945 ;
        RECT 60.715 24.775 61.005 24.945 ;
        RECT 61.175 24.775 61.465 24.945 ;
        RECT 61.635 24.775 61.925 24.945 ;
        RECT 62.095 24.775 62.385 24.945 ;
        RECT 62.555 24.775 62.845 24.945 ;
        RECT 63.015 24.775 63.305 24.945 ;
        RECT 63.475 24.775 63.765 24.945 ;
        RECT 63.935 24.775 64.225 24.945 ;
        RECT 64.395 24.775 64.685 24.945 ;
        RECT 64.855 24.775 65.145 24.945 ;
        RECT 65.315 24.775 65.605 24.945 ;
        RECT 65.775 24.775 66.065 24.945 ;
        RECT 66.235 24.775 66.525 24.945 ;
        RECT 66.695 24.775 66.985 24.945 ;
        RECT 67.155 24.775 67.445 24.945 ;
        RECT 67.615 24.775 67.905 24.945 ;
        RECT 68.075 24.775 68.365 24.945 ;
        RECT 68.535 24.775 68.825 24.945 ;
        RECT 68.995 24.775 69.285 24.945 ;
        RECT 69.455 24.775 69.745 24.945 ;
        RECT 69.915 24.775 70.205 24.945 ;
        RECT 70.375 24.775 70.665 24.945 ;
        RECT 70.835 24.775 71.125 24.945 ;
        RECT 71.295 24.775 71.585 24.945 ;
        RECT 71.755 24.775 72.045 24.945 ;
        RECT 72.215 24.775 72.505 24.945 ;
        RECT 72.675 24.775 72.965 24.945 ;
        RECT 73.135 24.775 73.425 24.945 ;
        RECT 73.595 24.775 73.885 24.945 ;
        RECT 74.055 24.775 74.345 24.945 ;
        RECT 74.515 24.775 74.805 24.945 ;
        RECT 74.975 24.775 75.265 24.945 ;
        RECT 75.435 24.775 75.725 24.945 ;
        RECT 75.895 24.775 76.185 24.945 ;
        RECT 76.355 24.775 76.645 24.945 ;
        RECT 76.815 24.775 77.105 24.945 ;
        RECT 77.275 24.775 77.565 24.945 ;
        RECT 77.735 24.775 78.025 24.945 ;
        RECT 78.195 24.775 78.485 24.945 ;
        RECT 78.655 24.775 78.945 24.945 ;
        RECT 79.115 24.775 79.405 24.945 ;
        RECT 79.575 24.775 79.865 24.945 ;
        RECT 80.035 24.775 80.325 24.945 ;
        RECT 80.495 24.775 80.785 24.945 ;
        RECT 80.955 24.775 81.245 24.945 ;
        RECT 81.415 24.775 81.705 24.945 ;
        RECT 81.875 24.775 82.165 24.945 ;
        RECT 82.335 24.775 82.625 24.945 ;
        RECT 82.795 24.775 83.085 24.945 ;
        RECT 83.255 24.775 83.545 24.945 ;
        RECT 83.715 24.775 84.005 24.945 ;
        RECT 84.175 24.775 84.465 24.945 ;
        RECT 84.635 24.775 84.925 24.945 ;
        RECT 85.095 24.775 85.385 24.945 ;
        RECT 85.555 24.775 85.845 24.945 ;
        RECT 86.015 24.775 86.305 24.945 ;
        RECT 86.475 24.775 86.765 24.945 ;
        RECT 86.935 24.775 87.225 24.945 ;
        RECT 87.395 24.775 87.685 24.945 ;
        RECT 87.855 24.775 88.145 24.945 ;
        RECT 88.315 24.775 88.605 24.945 ;
        RECT 88.775 24.775 89.065 24.945 ;
        RECT 89.235 24.775 89.525 24.945 ;
        RECT 89.695 24.775 89.985 24.945 ;
        RECT 90.155 24.775 90.445 24.945 ;
        RECT 90.615 24.775 90.905 24.945 ;
        RECT 91.075 24.775 91.365 24.945 ;
        RECT 91.535 24.775 91.825 24.945 ;
        RECT 91.995 24.775 92.285 24.945 ;
        RECT 92.455 24.775 92.745 24.945 ;
        RECT 92.915 24.775 93.205 24.945 ;
        RECT 93.375 24.775 93.665 24.945 ;
        RECT 93.835 24.775 94.125 24.945 ;
        RECT 94.295 24.775 94.585 24.945 ;
        RECT 94.755 24.775 95.045 24.945 ;
        RECT 95.215 24.775 95.505 24.945 ;
        RECT 95.675 24.775 95.965 24.945 ;
        RECT 96.135 24.775 96.425 24.945 ;
        RECT 96.595 24.775 96.885 24.945 ;
        RECT 97.055 24.775 97.345 24.945 ;
        RECT 97.515 24.775 97.805 24.945 ;
        RECT 97.975 24.775 98.265 24.945 ;
        RECT 98.435 24.775 98.725 24.945 ;
        RECT 98.895 24.775 99.185 24.945 ;
        RECT 99.355 24.775 99.645 24.945 ;
        RECT 99.815 24.775 99.960 24.945 ;
        RECT 16.785 24.025 17.995 24.775 ;
        RECT 16.785 23.485 17.305 24.025 ;
        RECT 18.165 24.005 23.510 24.775 ;
        RECT 23.685 24.005 29.030 24.775 ;
        RECT 29.205 24.005 30.875 24.775 ;
        RECT 31.045 24.050 31.335 24.775 ;
        RECT 31.505 24.005 36.850 24.775 ;
        RECT 37.025 24.005 42.370 24.775 ;
        RECT 42.545 24.005 47.890 24.775 ;
        RECT 48.065 24.005 53.410 24.775 ;
        RECT 53.585 24.005 58.930 24.775 ;
        RECT 59.105 24.050 59.395 24.775 ;
        RECT 59.565 24.005 64.910 24.775 ;
        RECT 65.085 24.005 70.430 24.775 ;
        RECT 70.605 24.005 72.275 24.775 ;
        RECT 72.915 24.245 73.245 24.605 ;
        RECT 73.775 24.415 74.105 24.775 ;
        RECT 74.710 24.415 75.040 24.775 ;
      LAYER li1 ;
        RECT 74.350 24.245 74.540 24.345 ;
        RECT 75.210 24.245 75.400 24.605 ;
      LAYER li1 ;
        RECT 75.570 24.415 75.900 24.775 ;
        RECT 72.915 24.055 74.180 24.245 ;
        RECT 17.475 23.315 17.995 23.855 ;
        RECT 18.165 23.485 20.745 24.005 ;
        RECT 20.915 23.315 23.510 23.835 ;
        RECT 23.685 23.485 26.265 24.005 ;
        RECT 26.435 23.315 29.030 23.835 ;
        RECT 29.205 23.485 29.955 24.005 ;
        RECT 30.125 23.315 30.875 23.835 ;
        RECT 31.505 23.485 34.085 24.005 ;
        RECT 16.785 22.225 17.995 23.315 ;
        RECT 18.165 22.225 23.510 23.315 ;
        RECT 23.685 22.225 29.030 23.315 ;
        RECT 29.205 22.225 30.875 23.315 ;
        RECT 31.045 22.225 31.335 23.390 ;
        RECT 34.255 23.315 36.850 23.835 ;
        RECT 37.025 23.485 39.605 24.005 ;
        RECT 39.775 23.315 42.370 23.835 ;
        RECT 42.545 23.485 45.125 24.005 ;
        RECT 45.295 23.315 47.890 23.835 ;
        RECT 48.065 23.485 50.645 24.005 ;
        RECT 50.815 23.315 53.410 23.835 ;
        RECT 53.585 23.485 56.165 24.005 ;
        RECT 56.335 23.315 58.930 23.835 ;
        RECT 59.565 23.485 62.145 24.005 ;
        RECT 31.505 22.225 36.850 23.315 ;
        RECT 37.025 22.225 42.370 23.315 ;
        RECT 42.545 22.225 47.890 23.315 ;
        RECT 48.065 22.225 53.410 23.315 ;
        RECT 53.585 22.225 58.930 23.315 ;
        RECT 59.105 22.225 59.395 23.390 ;
        RECT 62.315 23.315 64.910 23.835 ;
        RECT 65.085 23.485 67.665 24.005 ;
        RECT 67.835 23.315 70.430 23.835 ;
        RECT 70.605 23.485 71.355 24.005 ;
        RECT 71.525 23.315 72.275 23.835 ;
        RECT 59.565 22.225 64.910 23.315 ;
        RECT 65.085 22.225 70.430 23.315 ;
        RECT 70.605 22.225 72.275 23.315 ;
      LAYER li1 ;
        RECT 72.945 23.245 73.255 23.865 ;
      LAYER li1 ;
        RECT 73.970 23.840 74.180 24.055 ;
      LAYER li1 ;
        RECT 74.350 24.015 75.955 24.245 ;
      LAYER li1 ;
        RECT 73.970 23.505 75.505 23.840 ;
        RECT 73.970 23.280 74.180 23.505 ;
      LAYER li1 ;
        RECT 75.675 23.325 75.955 24.015 ;
      LAYER li1 ;
        RECT 76.125 24.005 81.470 24.775 ;
        RECT 81.645 24.005 86.990 24.775 ;
        RECT 87.165 24.050 87.455 24.775 ;
        RECT 87.625 24.005 92.970 24.775 ;
        RECT 93.145 24.005 98.490 24.775 ;
        RECT 98.665 24.025 99.875 24.775 ;
        RECT 76.125 23.485 78.705 24.005 ;
        RECT 73.425 23.110 74.180 23.280 ;
        RECT 72.915 22.225 73.245 22.980 ;
        RECT 73.425 22.395 73.605 23.110 ;
      LAYER li1 ;
        RECT 74.350 23.100 75.955 23.325 ;
      LAYER li1 ;
        RECT 78.875 23.315 81.470 23.835 ;
        RECT 81.645 23.485 84.225 24.005 ;
        RECT 84.395 23.315 86.990 23.835 ;
        RECT 87.625 23.485 90.205 24.005 ;
        RECT 73.810 22.225 74.140 22.925 ;
      LAYER li1 ;
        RECT 74.350 22.735 74.540 23.100 ;
        RECT 75.210 23.095 75.955 23.100 ;
        RECT 74.345 22.565 74.540 22.735 ;
        RECT 74.350 22.395 74.540 22.565 ;
      LAYER li1 ;
        RECT 74.710 22.225 75.040 22.925 ;
      LAYER li1 ;
        RECT 75.210 22.395 75.400 23.095 ;
      LAYER li1 ;
        RECT 75.570 22.225 75.900 22.925 ;
        RECT 76.125 22.225 81.470 23.315 ;
        RECT 81.645 22.225 86.990 23.315 ;
        RECT 87.165 22.225 87.455 23.390 ;
        RECT 90.375 23.315 92.970 23.835 ;
        RECT 93.145 23.485 95.725 24.005 ;
        RECT 95.895 23.315 98.490 23.835 ;
        RECT 87.625 22.225 92.970 23.315 ;
        RECT 93.145 22.225 98.490 23.315 ;
        RECT 98.665 23.315 99.185 23.855 ;
        RECT 99.355 23.485 99.875 24.025 ;
        RECT 98.665 22.225 99.875 23.315 ;
        RECT 16.700 22.055 16.845 22.225 ;
        RECT 17.015 22.055 17.305 22.225 ;
        RECT 17.475 22.055 17.765 22.225 ;
        RECT 17.935 22.055 18.225 22.225 ;
        RECT 18.395 22.055 18.685 22.225 ;
        RECT 18.855 22.055 19.145 22.225 ;
        RECT 19.315 22.055 19.605 22.225 ;
        RECT 19.775 22.055 20.065 22.225 ;
        RECT 20.235 22.055 20.525 22.225 ;
        RECT 20.695 22.055 20.985 22.225 ;
        RECT 21.155 22.055 21.445 22.225 ;
        RECT 21.615 22.055 21.905 22.225 ;
        RECT 22.075 22.055 22.365 22.225 ;
        RECT 22.535 22.055 22.825 22.225 ;
        RECT 22.995 22.055 23.285 22.225 ;
        RECT 23.455 22.055 23.745 22.225 ;
        RECT 23.915 22.055 24.205 22.225 ;
        RECT 24.375 22.055 24.665 22.225 ;
        RECT 24.835 22.055 25.125 22.225 ;
        RECT 25.295 22.055 25.585 22.225 ;
        RECT 25.755 22.055 26.045 22.225 ;
        RECT 26.215 22.055 26.505 22.225 ;
        RECT 26.675 22.055 26.965 22.225 ;
        RECT 27.135 22.055 27.425 22.225 ;
        RECT 27.595 22.055 27.885 22.225 ;
        RECT 28.055 22.055 28.345 22.225 ;
        RECT 28.515 22.055 28.805 22.225 ;
        RECT 28.975 22.055 29.265 22.225 ;
        RECT 29.435 22.055 29.725 22.225 ;
        RECT 29.895 22.055 30.185 22.225 ;
        RECT 30.355 22.055 30.645 22.225 ;
        RECT 30.815 22.055 31.105 22.225 ;
        RECT 31.275 22.055 31.565 22.225 ;
        RECT 31.735 22.055 32.025 22.225 ;
        RECT 32.195 22.055 32.485 22.225 ;
        RECT 32.655 22.055 32.945 22.225 ;
        RECT 33.115 22.055 33.405 22.225 ;
        RECT 33.575 22.055 33.865 22.225 ;
        RECT 34.035 22.055 34.325 22.225 ;
        RECT 34.495 22.055 34.785 22.225 ;
        RECT 34.955 22.055 35.245 22.225 ;
        RECT 35.415 22.055 35.705 22.225 ;
        RECT 35.875 22.055 36.165 22.225 ;
        RECT 36.335 22.055 36.625 22.225 ;
        RECT 36.795 22.055 37.085 22.225 ;
        RECT 37.255 22.055 37.545 22.225 ;
        RECT 37.715 22.055 38.005 22.225 ;
        RECT 38.175 22.055 38.465 22.225 ;
        RECT 38.635 22.055 38.925 22.225 ;
        RECT 39.095 22.055 39.385 22.225 ;
        RECT 39.555 22.055 39.845 22.225 ;
        RECT 40.015 22.055 40.305 22.225 ;
        RECT 40.475 22.055 40.765 22.225 ;
        RECT 40.935 22.055 41.225 22.225 ;
        RECT 41.395 22.055 41.685 22.225 ;
        RECT 41.855 22.055 42.145 22.225 ;
        RECT 42.315 22.055 42.605 22.225 ;
        RECT 42.775 22.055 43.065 22.225 ;
        RECT 43.235 22.055 43.525 22.225 ;
        RECT 43.695 22.055 43.985 22.225 ;
        RECT 44.155 22.055 44.445 22.225 ;
        RECT 44.615 22.055 44.905 22.225 ;
        RECT 45.075 22.055 45.365 22.225 ;
        RECT 45.535 22.055 45.825 22.225 ;
        RECT 45.995 22.055 46.285 22.225 ;
        RECT 46.455 22.055 46.745 22.225 ;
        RECT 46.915 22.055 47.205 22.225 ;
        RECT 47.375 22.055 47.665 22.225 ;
        RECT 47.835 22.055 48.125 22.225 ;
        RECT 48.295 22.055 48.585 22.225 ;
        RECT 48.755 22.055 49.045 22.225 ;
        RECT 49.215 22.055 49.505 22.225 ;
        RECT 49.675 22.055 49.965 22.225 ;
        RECT 50.135 22.055 50.425 22.225 ;
        RECT 50.595 22.055 50.885 22.225 ;
        RECT 51.055 22.055 51.345 22.225 ;
        RECT 51.515 22.055 51.805 22.225 ;
        RECT 51.975 22.055 52.265 22.225 ;
        RECT 52.435 22.055 52.725 22.225 ;
        RECT 52.895 22.055 53.185 22.225 ;
        RECT 53.355 22.055 53.645 22.225 ;
        RECT 53.815 22.055 54.105 22.225 ;
        RECT 54.275 22.055 54.565 22.225 ;
        RECT 54.735 22.055 55.025 22.225 ;
        RECT 55.195 22.055 55.485 22.225 ;
        RECT 55.655 22.055 55.945 22.225 ;
        RECT 56.115 22.055 56.405 22.225 ;
        RECT 56.575 22.055 56.865 22.225 ;
        RECT 57.035 22.055 57.325 22.225 ;
        RECT 57.495 22.055 57.785 22.225 ;
        RECT 57.955 22.055 58.245 22.225 ;
        RECT 58.415 22.055 58.705 22.225 ;
        RECT 58.875 22.055 59.165 22.225 ;
        RECT 59.335 22.055 59.625 22.225 ;
        RECT 59.795 22.055 60.085 22.225 ;
        RECT 60.255 22.055 60.545 22.225 ;
        RECT 60.715 22.055 61.005 22.225 ;
        RECT 61.175 22.055 61.465 22.225 ;
        RECT 61.635 22.055 61.925 22.225 ;
        RECT 62.095 22.055 62.385 22.225 ;
        RECT 62.555 22.055 62.845 22.225 ;
        RECT 63.015 22.055 63.305 22.225 ;
        RECT 63.475 22.055 63.765 22.225 ;
        RECT 63.935 22.055 64.225 22.225 ;
        RECT 64.395 22.055 64.685 22.225 ;
        RECT 64.855 22.055 65.145 22.225 ;
        RECT 65.315 22.055 65.605 22.225 ;
        RECT 65.775 22.055 66.065 22.225 ;
        RECT 66.235 22.055 66.525 22.225 ;
        RECT 66.695 22.055 66.985 22.225 ;
        RECT 67.155 22.055 67.445 22.225 ;
        RECT 67.615 22.055 67.905 22.225 ;
        RECT 68.075 22.055 68.365 22.225 ;
        RECT 68.535 22.055 68.825 22.225 ;
        RECT 68.995 22.055 69.285 22.225 ;
        RECT 69.455 22.055 69.745 22.225 ;
        RECT 69.915 22.055 70.205 22.225 ;
        RECT 70.375 22.055 70.665 22.225 ;
        RECT 70.835 22.055 71.125 22.225 ;
        RECT 71.295 22.055 71.585 22.225 ;
        RECT 71.755 22.055 72.045 22.225 ;
        RECT 72.215 22.055 72.505 22.225 ;
        RECT 72.675 22.055 72.965 22.225 ;
        RECT 73.135 22.055 73.425 22.225 ;
        RECT 73.595 22.055 73.885 22.225 ;
        RECT 74.055 22.055 74.345 22.225 ;
        RECT 74.515 22.055 74.805 22.225 ;
        RECT 74.975 22.055 75.265 22.225 ;
        RECT 75.435 22.055 75.725 22.225 ;
        RECT 75.895 22.055 76.185 22.225 ;
        RECT 76.355 22.055 76.645 22.225 ;
        RECT 76.815 22.055 77.105 22.225 ;
        RECT 77.275 22.055 77.565 22.225 ;
        RECT 77.735 22.055 78.025 22.225 ;
        RECT 78.195 22.055 78.485 22.225 ;
        RECT 78.655 22.055 78.945 22.225 ;
        RECT 79.115 22.055 79.405 22.225 ;
        RECT 79.575 22.055 79.865 22.225 ;
        RECT 80.035 22.055 80.325 22.225 ;
        RECT 80.495 22.055 80.785 22.225 ;
        RECT 80.955 22.055 81.245 22.225 ;
        RECT 81.415 22.055 81.705 22.225 ;
        RECT 81.875 22.055 82.165 22.225 ;
        RECT 82.335 22.055 82.625 22.225 ;
        RECT 82.795 22.055 83.085 22.225 ;
        RECT 83.255 22.055 83.545 22.225 ;
        RECT 83.715 22.055 84.005 22.225 ;
        RECT 84.175 22.055 84.465 22.225 ;
        RECT 84.635 22.055 84.925 22.225 ;
        RECT 85.095 22.055 85.385 22.225 ;
        RECT 85.555 22.055 85.845 22.225 ;
        RECT 86.015 22.055 86.305 22.225 ;
        RECT 86.475 22.055 86.765 22.225 ;
        RECT 86.935 22.055 87.225 22.225 ;
        RECT 87.395 22.055 87.685 22.225 ;
        RECT 87.855 22.055 88.145 22.225 ;
        RECT 88.315 22.055 88.605 22.225 ;
        RECT 88.775 22.055 89.065 22.225 ;
        RECT 89.235 22.055 89.525 22.225 ;
        RECT 89.695 22.055 89.985 22.225 ;
        RECT 90.155 22.055 90.445 22.225 ;
        RECT 90.615 22.055 90.905 22.225 ;
        RECT 91.075 22.055 91.365 22.225 ;
        RECT 91.535 22.055 91.825 22.225 ;
        RECT 91.995 22.055 92.285 22.225 ;
        RECT 92.455 22.055 92.745 22.225 ;
        RECT 92.915 22.055 93.205 22.225 ;
        RECT 93.375 22.055 93.665 22.225 ;
        RECT 93.835 22.055 94.125 22.225 ;
        RECT 94.295 22.055 94.585 22.225 ;
        RECT 94.755 22.055 95.045 22.225 ;
        RECT 95.215 22.055 95.505 22.225 ;
        RECT 95.675 22.055 95.965 22.225 ;
        RECT 96.135 22.055 96.425 22.225 ;
        RECT 96.595 22.055 96.885 22.225 ;
        RECT 97.055 22.055 97.345 22.225 ;
        RECT 97.515 22.055 97.805 22.225 ;
        RECT 97.975 22.055 98.265 22.225 ;
        RECT 98.435 22.055 98.725 22.225 ;
        RECT 98.895 22.055 99.185 22.225 ;
        RECT 99.355 22.055 99.645 22.225 ;
        RECT 99.815 22.055 99.960 22.225 ;
        RECT 16.785 20.965 17.995 22.055 ;
        RECT 18.165 20.965 19.375 22.055 ;
        RECT 19.735 21.330 20.065 22.055 ;
        RECT 16.785 20.255 17.305 20.795 ;
        RECT 17.475 20.425 17.995 20.965 ;
        RECT 18.165 20.255 18.685 20.795 ;
        RECT 18.855 20.425 19.375 20.965 ;
        RECT 16.785 19.505 17.995 20.255 ;
        RECT 18.165 19.505 19.375 20.255 ;
      LAYER li1 ;
        RECT 19.545 19.675 20.065 21.160 ;
      LAYER li1 ;
        RECT 20.925 20.965 26.270 22.055 ;
        RECT 26.445 20.965 31.790 22.055 ;
        RECT 31.965 20.965 37.310 22.055 ;
        RECT 37.485 20.965 42.830 22.055 ;
        RECT 43.005 20.965 44.675 22.055 ;
        RECT 20.925 20.275 23.505 20.795 ;
        RECT 23.675 20.445 26.270 20.965 ;
        RECT 26.445 20.275 29.025 20.795 ;
        RECT 29.195 20.445 31.790 20.965 ;
        RECT 31.965 20.275 34.545 20.795 ;
        RECT 34.715 20.445 37.310 20.965 ;
        RECT 37.485 20.275 40.065 20.795 ;
        RECT 40.235 20.445 42.830 20.965 ;
        RECT 43.005 20.275 43.755 20.795 ;
        RECT 43.925 20.445 44.675 20.965 ;
        RECT 44.845 20.890 45.135 22.055 ;
        RECT 45.305 20.965 50.650 22.055 ;
        RECT 50.825 20.965 53.415 22.055 ;
        RECT 54.135 21.385 54.305 21.885 ;
        RECT 54.475 21.555 54.805 22.055 ;
        RECT 54.135 21.215 54.800 21.385 ;
        RECT 45.305 20.275 47.885 20.795 ;
        RECT 48.055 20.445 50.650 20.965 ;
        RECT 50.825 20.275 52.035 20.795 ;
        RECT 52.205 20.445 53.415 20.965 ;
      LAYER li1 ;
        RECT 54.050 20.395 54.400 21.045 ;
      LAYER li1 ;
        RECT 20.235 19.505 20.575 20.165 ;
        RECT 20.925 19.505 26.270 20.275 ;
        RECT 26.445 19.505 31.790 20.275 ;
        RECT 31.965 19.505 37.310 20.275 ;
        RECT 37.485 19.505 42.830 20.275 ;
        RECT 43.005 19.505 44.675 20.275 ;
        RECT 44.845 19.505 45.135 20.230 ;
        RECT 45.305 19.505 50.650 20.275 ;
        RECT 50.825 19.505 53.415 20.275 ;
        RECT 54.570 20.225 54.800 21.215 ;
        RECT 54.135 20.055 54.800 20.225 ;
        RECT 54.135 19.765 54.305 20.055 ;
        RECT 54.475 19.505 54.805 19.885 ;
        RECT 54.975 19.765 55.200 21.885 ;
        RECT 55.400 21.595 55.665 22.055 ;
        RECT 55.850 21.485 56.085 21.860 ;
        RECT 56.330 21.610 57.400 21.780 ;
      LAYER li1 ;
        RECT 55.400 20.485 55.680 21.085 ;
      LAYER li1 ;
        RECT 55.415 19.505 55.665 19.965 ;
        RECT 55.850 19.955 56.020 21.485 ;
        RECT 56.190 20.455 56.430 21.325 ;
        RECT 56.620 21.075 57.060 21.430 ;
        RECT 57.230 20.995 57.400 21.610 ;
        RECT 57.570 21.255 57.740 22.055 ;
        RECT 57.910 21.555 58.160 21.885 ;
        RECT 58.385 21.585 59.270 21.755 ;
        RECT 57.230 20.905 57.740 20.995 ;
        RECT 56.940 20.735 57.740 20.905 ;
        RECT 56.190 20.125 56.770 20.455 ;
        RECT 56.940 19.955 57.110 20.735 ;
        RECT 57.570 20.665 57.740 20.735 ;
        RECT 57.280 20.485 57.450 20.515 ;
        RECT 57.910 20.485 58.080 21.555 ;
        RECT 58.250 20.665 58.440 21.385 ;
        RECT 58.610 20.995 58.930 21.325 ;
        RECT 57.280 20.185 58.080 20.485 ;
        RECT 58.610 20.455 58.800 20.995 ;
        RECT 55.850 19.785 56.180 19.955 ;
        RECT 56.360 19.785 57.110 19.955 ;
        RECT 57.360 19.505 57.730 20.005 ;
        RECT 57.910 19.955 58.080 20.185 ;
        RECT 58.250 20.125 58.800 20.455 ;
        RECT 59.100 20.665 59.270 21.585 ;
        RECT 59.450 21.555 59.665 22.055 ;
        RECT 60.130 21.250 60.300 21.875 ;
        RECT 60.585 21.275 60.765 22.055 ;
        RECT 59.440 21.090 60.300 21.250 ;
        RECT 61.460 21.225 61.630 22.055 ;
        RECT 62.300 21.225 62.470 22.055 ;
        RECT 59.440 20.920 60.550 21.090 ;
        RECT 62.785 20.965 68.130 22.055 ;
        RECT 68.305 20.965 71.815 22.055 ;
        RECT 60.380 20.665 60.550 20.920 ;
        RECT 59.100 20.495 60.190 20.665 ;
        RECT 60.380 20.495 62.200 20.665 ;
        RECT 59.100 19.955 59.270 20.495 ;
        RECT 60.380 20.325 60.550 20.495 ;
        RECT 60.050 20.155 60.550 20.325 ;
        RECT 62.785 20.275 65.365 20.795 ;
        RECT 65.535 20.445 68.130 20.965 ;
        RECT 68.305 20.275 69.955 20.795 ;
        RECT 70.125 20.445 71.815 20.965 ;
        RECT 72.905 20.890 73.195 22.055 ;
        RECT 73.455 21.385 73.625 21.885 ;
        RECT 73.795 21.555 74.125 22.055 ;
        RECT 73.455 21.215 74.120 21.385 ;
      LAYER li1 ;
        RECT 73.370 20.395 73.720 21.045 ;
      LAYER li1 ;
        RECT 57.910 19.785 58.370 19.955 ;
        RECT 58.600 19.785 59.270 19.955 ;
        RECT 59.585 19.505 59.755 20.035 ;
        RECT 60.050 19.715 60.410 20.155 ;
        RECT 60.585 19.505 60.755 19.985 ;
        RECT 61.455 19.505 61.625 19.980 ;
        RECT 62.305 19.505 62.475 19.980 ;
        RECT 62.785 19.505 68.130 20.275 ;
        RECT 68.305 19.505 71.815 20.275 ;
        RECT 72.905 19.505 73.195 20.230 ;
        RECT 73.890 20.225 74.120 21.215 ;
        RECT 73.455 20.055 74.120 20.225 ;
        RECT 73.455 19.765 73.625 20.055 ;
        RECT 73.795 19.505 74.125 19.885 ;
        RECT 74.295 19.765 74.520 21.885 ;
        RECT 74.720 21.595 74.985 22.055 ;
        RECT 75.170 21.485 75.405 21.860 ;
        RECT 75.650 21.610 76.720 21.780 ;
      LAYER li1 ;
        RECT 74.720 20.485 75.000 21.085 ;
      LAYER li1 ;
        RECT 74.735 19.505 74.985 19.965 ;
        RECT 75.170 19.955 75.340 21.485 ;
        RECT 75.510 20.455 75.750 21.325 ;
        RECT 75.940 21.075 76.380 21.430 ;
        RECT 76.550 20.995 76.720 21.610 ;
        RECT 76.890 21.255 77.060 22.055 ;
        RECT 77.230 21.555 77.480 21.885 ;
        RECT 77.705 21.585 78.590 21.755 ;
        RECT 76.550 20.905 77.060 20.995 ;
        RECT 76.260 20.735 77.060 20.905 ;
        RECT 75.510 20.125 76.090 20.455 ;
        RECT 76.260 19.955 76.430 20.735 ;
        RECT 76.890 20.665 77.060 20.735 ;
        RECT 76.600 20.485 76.770 20.515 ;
        RECT 77.230 20.485 77.400 21.555 ;
        RECT 77.570 20.665 77.760 21.385 ;
        RECT 77.930 20.995 78.250 21.325 ;
        RECT 76.600 20.185 77.400 20.485 ;
        RECT 77.930 20.455 78.120 20.995 ;
        RECT 75.170 19.785 75.500 19.955 ;
        RECT 75.680 19.785 76.430 19.955 ;
        RECT 76.680 19.505 77.050 20.005 ;
        RECT 77.230 19.955 77.400 20.185 ;
        RECT 77.570 20.125 78.120 20.455 ;
        RECT 78.420 20.665 78.590 21.585 ;
        RECT 78.770 21.555 78.985 22.055 ;
        RECT 79.450 21.250 79.620 21.875 ;
        RECT 79.905 21.275 80.085 22.055 ;
        RECT 78.760 21.090 79.620 21.250 ;
        RECT 80.780 21.225 80.950 22.055 ;
        RECT 81.620 21.225 81.790 22.055 ;
        RECT 78.760 20.920 79.870 21.090 ;
        RECT 82.105 20.965 87.450 22.055 ;
        RECT 87.625 20.965 92.970 22.055 ;
        RECT 93.145 20.965 98.490 22.055 ;
        RECT 79.700 20.665 79.870 20.920 ;
        RECT 78.420 20.495 79.510 20.665 ;
        RECT 79.700 20.495 81.520 20.665 ;
        RECT 78.420 19.955 78.590 20.495 ;
        RECT 79.700 20.325 79.870 20.495 ;
        RECT 79.370 20.155 79.870 20.325 ;
        RECT 82.105 20.275 84.685 20.795 ;
        RECT 84.855 20.445 87.450 20.965 ;
        RECT 87.625 20.275 90.205 20.795 ;
        RECT 90.375 20.445 92.970 20.965 ;
        RECT 93.145 20.275 95.725 20.795 ;
        RECT 95.895 20.445 98.490 20.965 ;
        RECT 98.665 20.965 99.875 22.055 ;
        RECT 98.665 20.425 99.185 20.965 ;
        RECT 77.230 19.785 77.690 19.955 ;
        RECT 77.920 19.785 78.590 19.955 ;
        RECT 78.905 19.505 79.075 20.035 ;
        RECT 79.370 19.715 79.730 20.155 ;
        RECT 79.905 19.505 80.075 19.985 ;
        RECT 80.775 19.505 80.945 19.980 ;
        RECT 81.625 19.505 81.795 19.980 ;
        RECT 82.105 19.505 87.450 20.275 ;
        RECT 87.625 19.505 92.970 20.275 ;
        RECT 93.145 19.505 98.490 20.275 ;
        RECT 99.355 20.255 99.875 20.795 ;
        RECT 98.665 19.505 99.875 20.255 ;
        RECT 16.700 19.335 16.845 19.505 ;
        RECT 17.015 19.335 17.305 19.505 ;
        RECT 17.475 19.335 17.765 19.505 ;
        RECT 17.935 19.335 18.225 19.505 ;
        RECT 18.395 19.335 18.685 19.505 ;
        RECT 18.855 19.335 19.145 19.505 ;
        RECT 19.315 19.335 19.605 19.505 ;
        RECT 19.775 19.335 20.065 19.505 ;
        RECT 20.235 19.335 20.525 19.505 ;
        RECT 20.695 19.335 20.985 19.505 ;
        RECT 21.155 19.335 21.445 19.505 ;
        RECT 21.615 19.335 21.905 19.505 ;
        RECT 22.075 19.335 22.365 19.505 ;
        RECT 22.535 19.335 22.825 19.505 ;
        RECT 22.995 19.335 23.285 19.505 ;
        RECT 23.455 19.335 23.745 19.505 ;
        RECT 23.915 19.335 24.205 19.505 ;
        RECT 24.375 19.335 24.665 19.505 ;
        RECT 24.835 19.335 25.125 19.505 ;
        RECT 25.295 19.335 25.585 19.505 ;
        RECT 25.755 19.335 26.045 19.505 ;
        RECT 26.215 19.335 26.505 19.505 ;
        RECT 26.675 19.335 26.965 19.505 ;
        RECT 27.135 19.335 27.425 19.505 ;
        RECT 27.595 19.335 27.885 19.505 ;
        RECT 28.055 19.335 28.345 19.505 ;
        RECT 28.515 19.335 28.805 19.505 ;
        RECT 28.975 19.335 29.265 19.505 ;
        RECT 29.435 19.335 29.725 19.505 ;
        RECT 29.895 19.335 30.185 19.505 ;
        RECT 30.355 19.335 30.645 19.505 ;
        RECT 30.815 19.335 31.105 19.505 ;
        RECT 31.275 19.335 31.565 19.505 ;
        RECT 31.735 19.335 32.025 19.505 ;
        RECT 32.195 19.335 32.485 19.505 ;
        RECT 32.655 19.335 32.945 19.505 ;
        RECT 33.115 19.335 33.405 19.505 ;
        RECT 33.575 19.335 33.865 19.505 ;
        RECT 34.035 19.335 34.325 19.505 ;
        RECT 34.495 19.335 34.785 19.505 ;
        RECT 34.955 19.335 35.245 19.505 ;
        RECT 35.415 19.335 35.705 19.505 ;
        RECT 35.875 19.335 36.165 19.505 ;
        RECT 36.335 19.335 36.625 19.505 ;
        RECT 36.795 19.335 37.085 19.505 ;
        RECT 37.255 19.335 37.545 19.505 ;
        RECT 37.715 19.335 38.005 19.505 ;
        RECT 38.175 19.335 38.465 19.505 ;
        RECT 38.635 19.335 38.925 19.505 ;
        RECT 39.095 19.335 39.385 19.505 ;
        RECT 39.555 19.335 39.845 19.505 ;
        RECT 40.015 19.335 40.305 19.505 ;
        RECT 40.475 19.335 40.765 19.505 ;
        RECT 40.935 19.335 41.225 19.505 ;
        RECT 41.395 19.335 41.685 19.505 ;
        RECT 41.855 19.335 42.145 19.505 ;
        RECT 42.315 19.335 42.605 19.505 ;
        RECT 42.775 19.335 43.065 19.505 ;
        RECT 43.235 19.335 43.525 19.505 ;
        RECT 43.695 19.335 43.985 19.505 ;
        RECT 44.155 19.335 44.445 19.505 ;
        RECT 44.615 19.335 44.905 19.505 ;
        RECT 45.075 19.335 45.365 19.505 ;
        RECT 45.535 19.335 45.825 19.505 ;
        RECT 45.995 19.335 46.285 19.505 ;
        RECT 46.455 19.335 46.745 19.505 ;
        RECT 46.915 19.335 47.205 19.505 ;
        RECT 47.375 19.335 47.665 19.505 ;
        RECT 47.835 19.335 48.125 19.505 ;
        RECT 48.295 19.335 48.585 19.505 ;
        RECT 48.755 19.335 49.045 19.505 ;
        RECT 49.215 19.335 49.505 19.505 ;
        RECT 49.675 19.335 49.965 19.505 ;
        RECT 50.135 19.335 50.425 19.505 ;
        RECT 50.595 19.335 50.885 19.505 ;
        RECT 51.055 19.335 51.345 19.505 ;
        RECT 51.515 19.335 51.805 19.505 ;
        RECT 51.975 19.335 52.265 19.505 ;
        RECT 52.435 19.335 52.725 19.505 ;
        RECT 52.895 19.335 53.185 19.505 ;
        RECT 53.355 19.335 53.645 19.505 ;
        RECT 53.815 19.335 54.105 19.505 ;
        RECT 54.275 19.335 54.565 19.505 ;
        RECT 54.735 19.335 55.025 19.505 ;
        RECT 55.195 19.335 55.485 19.505 ;
        RECT 55.655 19.335 55.945 19.505 ;
        RECT 56.115 19.335 56.405 19.505 ;
        RECT 56.575 19.335 56.865 19.505 ;
        RECT 57.035 19.335 57.325 19.505 ;
        RECT 57.495 19.335 57.785 19.505 ;
        RECT 57.955 19.335 58.245 19.505 ;
        RECT 58.415 19.335 58.705 19.505 ;
        RECT 58.875 19.335 59.165 19.505 ;
        RECT 59.335 19.335 59.625 19.505 ;
        RECT 59.795 19.335 60.085 19.505 ;
        RECT 60.255 19.335 60.545 19.505 ;
        RECT 60.715 19.335 61.005 19.505 ;
        RECT 61.175 19.335 61.465 19.505 ;
        RECT 61.635 19.335 61.925 19.505 ;
        RECT 62.095 19.335 62.385 19.505 ;
        RECT 62.555 19.335 62.845 19.505 ;
        RECT 63.015 19.335 63.305 19.505 ;
        RECT 63.475 19.335 63.765 19.505 ;
        RECT 63.935 19.335 64.225 19.505 ;
        RECT 64.395 19.335 64.685 19.505 ;
        RECT 64.855 19.335 65.145 19.505 ;
        RECT 65.315 19.335 65.605 19.505 ;
        RECT 65.775 19.335 66.065 19.505 ;
        RECT 66.235 19.335 66.525 19.505 ;
        RECT 66.695 19.335 66.985 19.505 ;
        RECT 67.155 19.335 67.445 19.505 ;
        RECT 67.615 19.335 67.905 19.505 ;
        RECT 68.075 19.335 68.365 19.505 ;
        RECT 68.535 19.335 68.825 19.505 ;
        RECT 68.995 19.335 69.285 19.505 ;
        RECT 69.455 19.335 69.745 19.505 ;
        RECT 69.915 19.335 70.205 19.505 ;
        RECT 70.375 19.335 70.665 19.505 ;
        RECT 70.835 19.335 71.125 19.505 ;
        RECT 71.295 19.335 71.585 19.505 ;
        RECT 71.755 19.335 72.045 19.505 ;
        RECT 72.215 19.335 72.505 19.505 ;
        RECT 72.675 19.335 72.965 19.505 ;
        RECT 73.135 19.335 73.425 19.505 ;
        RECT 73.595 19.335 73.885 19.505 ;
        RECT 74.055 19.335 74.345 19.505 ;
        RECT 74.515 19.335 74.805 19.505 ;
        RECT 74.975 19.335 75.265 19.505 ;
        RECT 75.435 19.335 75.725 19.505 ;
        RECT 75.895 19.335 76.185 19.505 ;
        RECT 76.355 19.335 76.645 19.505 ;
        RECT 76.815 19.335 77.105 19.505 ;
        RECT 77.275 19.335 77.565 19.505 ;
        RECT 77.735 19.335 78.025 19.505 ;
        RECT 78.195 19.335 78.485 19.505 ;
        RECT 78.655 19.335 78.945 19.505 ;
        RECT 79.115 19.335 79.405 19.505 ;
        RECT 79.575 19.335 79.865 19.505 ;
        RECT 80.035 19.335 80.325 19.505 ;
        RECT 80.495 19.335 80.785 19.505 ;
        RECT 80.955 19.335 81.245 19.505 ;
        RECT 81.415 19.335 81.705 19.505 ;
        RECT 81.875 19.335 82.165 19.505 ;
        RECT 82.335 19.335 82.625 19.505 ;
        RECT 82.795 19.335 83.085 19.505 ;
        RECT 83.255 19.335 83.545 19.505 ;
        RECT 83.715 19.335 84.005 19.505 ;
        RECT 84.175 19.335 84.465 19.505 ;
        RECT 84.635 19.335 84.925 19.505 ;
        RECT 85.095 19.335 85.385 19.505 ;
        RECT 85.555 19.335 85.845 19.505 ;
        RECT 86.015 19.335 86.305 19.505 ;
        RECT 86.475 19.335 86.765 19.505 ;
        RECT 86.935 19.335 87.225 19.505 ;
        RECT 87.395 19.335 87.685 19.505 ;
        RECT 87.855 19.335 88.145 19.505 ;
        RECT 88.315 19.335 88.605 19.505 ;
        RECT 88.775 19.335 89.065 19.505 ;
        RECT 89.235 19.335 89.525 19.505 ;
        RECT 89.695 19.335 89.985 19.505 ;
        RECT 90.155 19.335 90.445 19.505 ;
        RECT 90.615 19.335 90.905 19.505 ;
        RECT 91.075 19.335 91.365 19.505 ;
        RECT 91.535 19.335 91.825 19.505 ;
        RECT 91.995 19.335 92.285 19.505 ;
        RECT 92.455 19.335 92.745 19.505 ;
        RECT 92.915 19.335 93.205 19.505 ;
        RECT 93.375 19.335 93.665 19.505 ;
        RECT 93.835 19.335 94.125 19.505 ;
        RECT 94.295 19.335 94.585 19.505 ;
        RECT 94.755 19.335 95.045 19.505 ;
        RECT 95.215 19.335 95.505 19.505 ;
        RECT 95.675 19.335 95.965 19.505 ;
        RECT 96.135 19.335 96.425 19.505 ;
        RECT 96.595 19.335 96.885 19.505 ;
        RECT 97.055 19.335 97.345 19.505 ;
        RECT 97.515 19.335 97.805 19.505 ;
        RECT 97.975 19.335 98.265 19.505 ;
        RECT 98.435 19.335 98.725 19.505 ;
        RECT 98.895 19.335 99.185 19.505 ;
        RECT 99.355 19.335 99.645 19.505 ;
        RECT 99.815 19.335 99.960 19.505 ;
        RECT 16.785 18.585 17.995 19.335 ;
        RECT 16.785 18.045 17.305 18.585 ;
        RECT 18.165 18.565 23.510 19.335 ;
        RECT 23.685 18.565 29.030 19.335 ;
        RECT 29.205 18.565 30.875 19.335 ;
        RECT 31.045 18.610 31.335 19.335 ;
        RECT 17.475 17.875 17.995 18.415 ;
        RECT 18.165 18.045 20.745 18.565 ;
        RECT 20.915 17.875 23.510 18.395 ;
        RECT 23.685 18.045 26.265 18.565 ;
        RECT 26.435 17.875 29.030 18.395 ;
        RECT 29.205 18.045 29.955 18.565 ;
        RECT 30.125 17.875 30.875 18.395 ;
        RECT 16.785 16.785 17.995 17.875 ;
        RECT 18.165 16.785 23.510 17.875 ;
        RECT 23.685 16.785 29.030 17.875 ;
        RECT 29.205 16.785 30.875 17.875 ;
        RECT 31.045 16.785 31.335 17.950 ;
      LAYER li1 ;
        RECT 31.505 17.680 32.025 19.165 ;
      LAYER li1 ;
        RECT 32.195 18.675 32.535 19.335 ;
        RECT 32.885 18.565 38.230 19.335 ;
        RECT 38.405 18.565 43.750 19.335 ;
        RECT 43.925 18.585 45.135 19.335 ;
        RECT 45.305 18.610 45.595 19.335 ;
        RECT 32.885 18.045 35.465 18.565 ;
        RECT 35.635 17.875 38.230 18.395 ;
        RECT 38.405 18.045 40.985 18.565 ;
        RECT 41.155 17.875 43.750 18.395 ;
        RECT 43.925 18.045 44.445 18.585 ;
        RECT 45.765 18.565 48.355 19.335 ;
        RECT 44.615 17.875 45.135 18.415 ;
        RECT 45.765 18.045 46.975 18.565 ;
        RECT 31.695 16.785 32.025 17.510 ;
        RECT 32.885 16.785 38.230 17.875 ;
        RECT 38.405 16.785 43.750 17.875 ;
        RECT 43.925 16.785 45.135 17.875 ;
        RECT 45.305 16.785 45.595 17.950 ;
        RECT 47.145 17.875 48.355 18.395 ;
        RECT 45.765 16.785 48.355 17.875 ;
      LAYER li1 ;
        RECT 48.985 17.680 49.505 19.165 ;
      LAYER li1 ;
        RECT 49.675 18.675 50.015 19.335 ;
        RECT 50.365 18.565 55.710 19.335 ;
        RECT 55.885 18.565 59.395 19.335 ;
        RECT 59.565 18.610 59.855 19.335 ;
        RECT 60.035 18.805 60.365 19.165 ;
        RECT 60.895 18.975 61.225 19.335 ;
        RECT 61.830 18.975 62.160 19.335 ;
      LAYER li1 ;
        RECT 61.470 18.805 61.660 18.905 ;
        RECT 62.330 18.805 62.520 19.165 ;
      LAYER li1 ;
        RECT 62.690 18.975 63.020 19.335 ;
        RECT 60.035 18.615 61.300 18.805 ;
        RECT 50.365 18.045 52.945 18.565 ;
        RECT 53.115 17.875 55.710 18.395 ;
        RECT 55.885 18.045 57.535 18.565 ;
        RECT 57.705 17.875 59.395 18.395 ;
        RECT 49.175 16.785 49.505 17.510 ;
        RECT 50.365 16.785 55.710 17.875 ;
        RECT 55.885 16.785 59.395 17.875 ;
        RECT 59.565 16.785 59.855 17.950 ;
      LAYER li1 ;
        RECT 60.065 17.805 60.375 18.425 ;
      LAYER li1 ;
        RECT 61.090 18.400 61.300 18.615 ;
      LAYER li1 ;
        RECT 61.470 18.575 63.075 18.805 ;
      LAYER li1 ;
        RECT 61.090 18.065 62.625 18.400 ;
        RECT 61.090 17.840 61.300 18.065 ;
      LAYER li1 ;
        RECT 62.795 17.885 63.075 18.575 ;
      LAYER li1 ;
        RECT 63.245 18.565 68.590 19.335 ;
        RECT 68.765 18.565 72.275 19.335 ;
        RECT 72.445 18.585 73.655 19.335 ;
        RECT 73.825 18.610 74.115 19.335 ;
        RECT 63.245 18.045 65.825 18.565 ;
        RECT 60.545 17.670 61.300 17.840 ;
        RECT 60.035 16.785 60.365 17.540 ;
        RECT 60.545 16.955 60.725 17.670 ;
      LAYER li1 ;
        RECT 61.470 17.660 63.075 17.885 ;
      LAYER li1 ;
        RECT 65.995 17.875 68.590 18.395 ;
        RECT 68.765 18.045 70.415 18.565 ;
        RECT 70.585 17.875 72.275 18.395 ;
        RECT 72.445 18.045 72.965 18.585 ;
        RECT 74.285 18.565 79.630 19.335 ;
        RECT 79.805 18.565 85.150 19.335 ;
        RECT 85.325 18.565 87.915 19.335 ;
        RECT 88.085 18.610 88.375 19.335 ;
        RECT 73.135 17.875 73.655 18.415 ;
        RECT 74.285 18.045 76.865 18.565 ;
        RECT 60.930 16.785 61.260 17.485 ;
      LAYER li1 ;
        RECT 61.470 17.295 61.660 17.660 ;
        RECT 62.330 17.655 63.075 17.660 ;
        RECT 61.465 17.125 61.660 17.295 ;
        RECT 61.470 16.955 61.660 17.125 ;
      LAYER li1 ;
        RECT 61.830 16.785 62.160 17.485 ;
      LAYER li1 ;
        RECT 62.330 16.955 62.520 17.655 ;
      LAYER li1 ;
        RECT 62.690 16.785 63.020 17.485 ;
        RECT 63.245 16.785 68.590 17.875 ;
        RECT 68.765 16.785 72.275 17.875 ;
        RECT 72.445 16.785 73.655 17.875 ;
        RECT 73.825 16.785 74.115 17.950 ;
        RECT 77.035 17.875 79.630 18.395 ;
        RECT 79.805 18.045 82.385 18.565 ;
        RECT 82.555 17.875 85.150 18.395 ;
        RECT 85.325 18.045 86.535 18.565 ;
        RECT 86.705 17.875 87.915 18.395 ;
        RECT 74.285 16.785 79.630 17.875 ;
        RECT 79.805 16.785 85.150 17.875 ;
        RECT 85.325 16.785 87.915 17.875 ;
        RECT 88.085 16.785 88.375 17.950 ;
      LAYER li1 ;
        RECT 88.545 17.680 89.065 19.165 ;
      LAYER li1 ;
        RECT 89.235 18.675 89.575 19.335 ;
        RECT 89.925 18.565 93.435 19.335 ;
        RECT 89.925 18.045 91.575 18.565 ;
        RECT 91.745 17.875 93.435 18.395 ;
        RECT 88.735 16.785 89.065 17.510 ;
        RECT 89.925 16.785 93.435 17.875 ;
      LAYER li1 ;
        RECT 93.605 17.680 94.125 19.165 ;
      LAYER li1 ;
        RECT 94.295 18.675 94.635 19.335 ;
        RECT 94.985 18.565 98.495 19.335 ;
        RECT 98.665 18.585 99.875 19.335 ;
        RECT 94.985 18.045 96.635 18.565 ;
        RECT 96.805 17.875 98.495 18.395 ;
        RECT 93.795 16.785 94.125 17.510 ;
        RECT 94.985 16.785 98.495 17.875 ;
        RECT 98.665 17.875 99.185 18.415 ;
        RECT 99.355 18.045 99.875 18.585 ;
        RECT 98.665 16.785 99.875 17.875 ;
        RECT 16.700 16.615 16.845 16.785 ;
        RECT 17.015 16.615 17.305 16.785 ;
        RECT 17.475 16.615 17.765 16.785 ;
        RECT 17.935 16.615 18.225 16.785 ;
        RECT 18.395 16.615 18.685 16.785 ;
        RECT 18.855 16.615 19.145 16.785 ;
        RECT 19.315 16.615 19.605 16.785 ;
        RECT 19.775 16.615 20.065 16.785 ;
        RECT 20.235 16.615 20.525 16.785 ;
        RECT 20.695 16.615 20.985 16.785 ;
        RECT 21.155 16.615 21.445 16.785 ;
        RECT 21.615 16.615 21.905 16.785 ;
        RECT 22.075 16.615 22.365 16.785 ;
        RECT 22.535 16.615 22.825 16.785 ;
        RECT 22.995 16.615 23.285 16.785 ;
        RECT 23.455 16.615 23.745 16.785 ;
        RECT 23.915 16.615 24.205 16.785 ;
        RECT 24.375 16.615 24.665 16.785 ;
        RECT 24.835 16.615 25.125 16.785 ;
        RECT 25.295 16.615 25.585 16.785 ;
        RECT 25.755 16.615 26.045 16.785 ;
        RECT 26.215 16.615 26.505 16.785 ;
        RECT 26.675 16.615 26.965 16.785 ;
        RECT 27.135 16.615 27.425 16.785 ;
        RECT 27.595 16.615 27.885 16.785 ;
        RECT 28.055 16.615 28.345 16.785 ;
        RECT 28.515 16.615 28.805 16.785 ;
        RECT 28.975 16.615 29.265 16.785 ;
        RECT 29.435 16.615 29.725 16.785 ;
        RECT 29.895 16.615 30.185 16.785 ;
        RECT 30.355 16.615 30.645 16.785 ;
        RECT 30.815 16.615 31.105 16.785 ;
        RECT 31.275 16.615 31.565 16.785 ;
        RECT 31.735 16.615 32.025 16.785 ;
        RECT 32.195 16.615 32.485 16.785 ;
        RECT 32.655 16.615 32.945 16.785 ;
        RECT 33.115 16.615 33.405 16.785 ;
        RECT 33.575 16.615 33.865 16.785 ;
        RECT 34.035 16.615 34.325 16.785 ;
        RECT 34.495 16.615 34.785 16.785 ;
        RECT 34.955 16.615 35.245 16.785 ;
        RECT 35.415 16.615 35.705 16.785 ;
        RECT 35.875 16.615 36.165 16.785 ;
        RECT 36.335 16.615 36.625 16.785 ;
        RECT 36.795 16.615 37.085 16.785 ;
        RECT 37.255 16.615 37.545 16.785 ;
        RECT 37.715 16.615 38.005 16.785 ;
        RECT 38.175 16.615 38.465 16.785 ;
        RECT 38.635 16.615 38.925 16.785 ;
        RECT 39.095 16.615 39.385 16.785 ;
        RECT 39.555 16.615 39.845 16.785 ;
        RECT 40.015 16.615 40.305 16.785 ;
        RECT 40.475 16.615 40.765 16.785 ;
        RECT 40.935 16.615 41.225 16.785 ;
        RECT 41.395 16.615 41.685 16.785 ;
        RECT 41.855 16.615 42.145 16.785 ;
        RECT 42.315 16.615 42.605 16.785 ;
        RECT 42.775 16.615 43.065 16.785 ;
        RECT 43.235 16.615 43.525 16.785 ;
        RECT 43.695 16.615 43.985 16.785 ;
        RECT 44.155 16.615 44.445 16.785 ;
        RECT 44.615 16.615 44.905 16.785 ;
        RECT 45.075 16.615 45.365 16.785 ;
        RECT 45.535 16.615 45.825 16.785 ;
        RECT 45.995 16.615 46.285 16.785 ;
        RECT 46.455 16.615 46.745 16.785 ;
        RECT 46.915 16.615 47.205 16.785 ;
        RECT 47.375 16.615 47.665 16.785 ;
        RECT 47.835 16.615 48.125 16.785 ;
        RECT 48.295 16.615 48.585 16.785 ;
        RECT 48.755 16.615 49.045 16.785 ;
        RECT 49.215 16.615 49.505 16.785 ;
        RECT 49.675 16.615 49.965 16.785 ;
        RECT 50.135 16.615 50.425 16.785 ;
        RECT 50.595 16.615 50.885 16.785 ;
        RECT 51.055 16.615 51.345 16.785 ;
        RECT 51.515 16.615 51.805 16.785 ;
        RECT 51.975 16.615 52.265 16.785 ;
        RECT 52.435 16.615 52.725 16.785 ;
        RECT 52.895 16.615 53.185 16.785 ;
        RECT 53.355 16.615 53.645 16.785 ;
        RECT 53.815 16.615 54.105 16.785 ;
        RECT 54.275 16.615 54.565 16.785 ;
        RECT 54.735 16.615 55.025 16.785 ;
        RECT 55.195 16.615 55.485 16.785 ;
        RECT 55.655 16.615 55.945 16.785 ;
        RECT 56.115 16.615 56.405 16.785 ;
        RECT 56.575 16.615 56.865 16.785 ;
        RECT 57.035 16.615 57.325 16.785 ;
        RECT 57.495 16.615 57.785 16.785 ;
        RECT 57.955 16.615 58.245 16.785 ;
        RECT 58.415 16.615 58.705 16.785 ;
        RECT 58.875 16.615 59.165 16.785 ;
        RECT 59.335 16.615 59.625 16.785 ;
        RECT 59.795 16.615 60.085 16.785 ;
        RECT 60.255 16.615 60.545 16.785 ;
        RECT 60.715 16.615 61.005 16.785 ;
        RECT 61.175 16.615 61.465 16.785 ;
        RECT 61.635 16.615 61.925 16.785 ;
        RECT 62.095 16.615 62.385 16.785 ;
        RECT 62.555 16.615 62.845 16.785 ;
        RECT 63.015 16.615 63.305 16.785 ;
        RECT 63.475 16.615 63.765 16.785 ;
        RECT 63.935 16.615 64.225 16.785 ;
        RECT 64.395 16.615 64.685 16.785 ;
        RECT 64.855 16.615 65.145 16.785 ;
        RECT 65.315 16.615 65.605 16.785 ;
        RECT 65.775 16.615 66.065 16.785 ;
        RECT 66.235 16.615 66.525 16.785 ;
        RECT 66.695 16.615 66.985 16.785 ;
        RECT 67.155 16.615 67.445 16.785 ;
        RECT 67.615 16.615 67.905 16.785 ;
        RECT 68.075 16.615 68.365 16.785 ;
        RECT 68.535 16.615 68.825 16.785 ;
        RECT 68.995 16.615 69.285 16.785 ;
        RECT 69.455 16.615 69.745 16.785 ;
        RECT 69.915 16.615 70.205 16.785 ;
        RECT 70.375 16.615 70.665 16.785 ;
        RECT 70.835 16.615 71.125 16.785 ;
        RECT 71.295 16.615 71.585 16.785 ;
        RECT 71.755 16.615 72.045 16.785 ;
        RECT 72.215 16.615 72.505 16.785 ;
        RECT 72.675 16.615 72.965 16.785 ;
        RECT 73.135 16.615 73.425 16.785 ;
        RECT 73.595 16.615 73.885 16.785 ;
        RECT 74.055 16.615 74.345 16.785 ;
        RECT 74.515 16.615 74.805 16.785 ;
        RECT 74.975 16.615 75.265 16.785 ;
        RECT 75.435 16.615 75.725 16.785 ;
        RECT 75.895 16.615 76.185 16.785 ;
        RECT 76.355 16.615 76.645 16.785 ;
        RECT 76.815 16.615 77.105 16.785 ;
        RECT 77.275 16.615 77.565 16.785 ;
        RECT 77.735 16.615 78.025 16.785 ;
        RECT 78.195 16.615 78.485 16.785 ;
        RECT 78.655 16.615 78.945 16.785 ;
        RECT 79.115 16.615 79.405 16.785 ;
        RECT 79.575 16.615 79.865 16.785 ;
        RECT 80.035 16.615 80.325 16.785 ;
        RECT 80.495 16.615 80.785 16.785 ;
        RECT 80.955 16.615 81.245 16.785 ;
        RECT 81.415 16.615 81.705 16.785 ;
        RECT 81.875 16.615 82.165 16.785 ;
        RECT 82.335 16.615 82.625 16.785 ;
        RECT 82.795 16.615 83.085 16.785 ;
        RECT 83.255 16.615 83.545 16.785 ;
        RECT 83.715 16.615 84.005 16.785 ;
        RECT 84.175 16.615 84.465 16.785 ;
        RECT 84.635 16.615 84.925 16.785 ;
        RECT 85.095 16.615 85.385 16.785 ;
        RECT 85.555 16.615 85.845 16.785 ;
        RECT 86.015 16.615 86.305 16.785 ;
        RECT 86.475 16.615 86.765 16.785 ;
        RECT 86.935 16.615 87.225 16.785 ;
        RECT 87.395 16.615 87.685 16.785 ;
        RECT 87.855 16.615 88.145 16.785 ;
        RECT 88.315 16.615 88.605 16.785 ;
        RECT 88.775 16.615 89.065 16.785 ;
        RECT 89.235 16.615 89.525 16.785 ;
        RECT 89.695 16.615 89.985 16.785 ;
        RECT 90.155 16.615 90.445 16.785 ;
        RECT 90.615 16.615 90.905 16.785 ;
        RECT 91.075 16.615 91.365 16.785 ;
        RECT 91.535 16.615 91.825 16.785 ;
        RECT 91.995 16.615 92.285 16.785 ;
        RECT 92.455 16.615 92.745 16.785 ;
        RECT 92.915 16.615 93.205 16.785 ;
        RECT 93.375 16.615 93.665 16.785 ;
        RECT 93.835 16.615 94.125 16.785 ;
        RECT 94.295 16.615 94.585 16.785 ;
        RECT 94.755 16.615 95.045 16.785 ;
        RECT 95.215 16.615 95.505 16.785 ;
        RECT 95.675 16.615 95.965 16.785 ;
        RECT 96.135 16.615 96.425 16.785 ;
        RECT 96.595 16.615 96.885 16.785 ;
        RECT 97.055 16.615 97.345 16.785 ;
        RECT 97.515 16.615 97.805 16.785 ;
        RECT 97.975 16.615 98.265 16.785 ;
        RECT 98.435 16.615 98.725 16.785 ;
        RECT 98.895 16.615 99.185 16.785 ;
        RECT 99.355 16.615 99.645 16.785 ;
        RECT 99.815 16.615 99.960 16.785 ;
      LAYER mcon ;
        RECT 64.225 91.245 64.395 91.415 ;
        RECT 66.985 90.905 67.155 91.075 ;
        RECT 62.385 88.865 62.555 89.035 ;
        RECT 63.765 88.865 63.935 89.035 ;
        RECT 35.705 82.405 35.875 82.575 ;
        RECT 38.005 80.365 38.175 80.535 ;
        RECT 40.765 80.025 40.935 80.195 ;
        RECT 38.925 77.645 39.095 77.815 ;
        RECT 40.305 77.985 40.475 78.155 ;
        RECT 73.425 77.645 73.595 77.815 ;
        RECT 74.805 77.985 74.975 78.155 ;
        RECT 56.865 67.785 57.035 67.955 ;
        RECT 57.785 67.105 57.955 67.275 ;
        RECT 60.545 64.045 60.715 64.215 ;
        RECT 61.925 64.045 62.095 64.215 ;
        RECT 40.765 61.665 40.935 61.835 ;
        RECT 42.145 61.325 42.315 61.495 ;
        RECT 60.085 61.665 60.255 61.835 ;
        RECT 61.005 60.645 61.175 60.815 ;
        RECT 68.825 61.325 68.995 61.495 ;
        RECT 70.205 61.325 70.375 61.495 ;
        RECT 40.765 58.945 40.935 59.115 ;
        RECT 38.465 58.605 38.635 58.775 ;
        RECT 63.765 58.605 63.935 58.775 ;
        RECT 65.145 55.885 65.315 56.055 ;
        RECT 67.905 56.565 68.075 56.735 ;
        RECT 62.845 53.845 63.015 54.015 ;
        RECT 61.005 50.785 61.175 50.955 ;
        RECT 62.385 50.445 62.555 50.615 ;
        RECT 59.625 48.745 59.795 48.915 ;
        RECT 60.545 47.725 60.715 47.895 ;
        RECT 59.625 45.005 59.795 45.175 ;
        RECT 62.385 45.685 62.555 45.855 ;
        RECT 72.965 23.585 73.135 23.755 ;
        RECT 54.105 20.865 54.275 21.035 ;
        RECT 55.485 20.525 55.655 20.695 ;
        RECT 73.425 20.865 73.595 21.035 ;
        RECT 74.805 20.865 74.975 21.035 ;
        RECT 60.085 18.145 60.255 18.315 ;
      LAYER met1 ;
        RECT 64.150 91.400 64.470 91.460 ;
        RECT 63.955 91.260 64.470 91.400 ;
        RECT 64.150 91.200 64.470 91.260 ;
        RECT 63.690 91.060 64.010 91.120 ;
        RECT 66.925 91.060 67.215 91.105 ;
        RECT 63.690 90.920 67.215 91.060 ;
        RECT 63.690 90.860 64.010 90.920 ;
        RECT 66.925 90.875 67.215 90.920 ;
      LAYER met1 ;
        RECT 63.250 89.360 63.540 89.405 ;
        RECT 64.650 89.360 64.940 89.405 ;
        RECT 66.490 89.360 66.780 89.405 ;
        RECT 63.250 89.220 66.780 89.360 ;
        RECT 63.250 89.175 63.540 89.220 ;
        RECT 64.650 89.175 64.940 89.220 ;
        RECT 66.490 89.175 66.780 89.220 ;
      LAYER met1 ;
        RECT 59.550 89.020 59.870 89.080 ;
        RECT 62.325 89.020 62.615 89.065 ;
        RECT 63.690 89.020 64.010 89.080 ;
        RECT 59.550 88.880 62.615 89.020 ;
        RECT 63.495 88.880 64.010 89.020 ;
        RECT 59.550 88.820 59.870 88.880 ;
        RECT 62.325 88.835 62.615 88.880 ;
        RECT 63.690 88.820 64.010 88.880 ;
      LAYER met1 ;
        RECT 62.790 88.340 63.080 88.385 ;
        RECT 65.110 88.340 65.400 88.385 ;
        RECT 66.490 88.340 66.780 88.385 ;
        RECT 62.790 88.200 66.780 88.340 ;
        RECT 62.790 88.155 63.080 88.200 ;
        RECT 65.110 88.155 65.400 88.200 ;
        RECT 66.490 88.155 66.780 88.200 ;
      LAYER met1 ;
        RECT 35.645 82.560 35.935 82.605 ;
        RECT 37.930 82.560 38.250 82.620 ;
        RECT 35.645 82.420 38.250 82.560 ;
        RECT 35.645 82.375 35.935 82.420 ;
        RECT 37.930 82.360 38.250 82.420 ;
        RECT 37.930 80.520 38.250 80.580 ;
        RECT 37.735 80.380 38.250 80.520 ;
        RECT 37.930 80.320 38.250 80.380 ;
        RECT 40.230 80.180 40.550 80.240 ;
        RECT 40.705 80.180 40.995 80.225 ;
        RECT 40.230 80.040 40.995 80.180 ;
        RECT 40.230 79.980 40.550 80.040 ;
        RECT 40.705 79.995 40.995 80.040 ;
      LAYER met1 ;
        RECT 39.790 78.480 40.080 78.525 ;
        RECT 41.190 78.480 41.480 78.525 ;
        RECT 43.030 78.480 43.320 78.525 ;
        RECT 39.790 78.340 43.320 78.480 ;
        RECT 39.790 78.295 40.080 78.340 ;
        RECT 41.190 78.295 41.480 78.340 ;
        RECT 43.030 78.295 43.320 78.340 ;
        RECT 74.290 78.480 74.580 78.525 ;
        RECT 75.690 78.480 75.980 78.525 ;
        RECT 77.530 78.480 77.820 78.525 ;
        RECT 74.290 78.340 77.820 78.480 ;
        RECT 74.290 78.295 74.580 78.340 ;
        RECT 75.690 78.295 75.980 78.340 ;
        RECT 77.530 78.295 77.820 78.340 ;
      LAYER met1 ;
        RECT 40.230 78.140 40.550 78.200 ;
        RECT 40.035 78.000 40.550 78.140 ;
        RECT 40.230 77.940 40.550 78.000 ;
        RECT 63.690 78.140 64.010 78.200 ;
        RECT 74.745 78.140 75.035 78.185 ;
        RECT 63.690 78.000 75.035 78.140 ;
        RECT 63.690 77.940 64.010 78.000 ;
        RECT 74.745 77.955 75.035 78.000 ;
        RECT 38.865 77.800 39.155 77.845 ;
        RECT 40.690 77.800 41.010 77.860 ;
        RECT 38.865 77.660 41.010 77.800 ;
        RECT 38.865 77.615 39.155 77.660 ;
        RECT 40.690 77.600 41.010 77.660 ;
        RECT 73.365 77.615 73.655 77.845 ;
      LAYER met1 ;
        RECT 39.330 77.460 39.620 77.505 ;
        RECT 41.650 77.460 41.940 77.505 ;
        RECT 43.030 77.460 43.320 77.505 ;
        RECT 39.330 77.320 43.320 77.460 ;
        RECT 39.330 77.275 39.620 77.320 ;
        RECT 41.650 77.275 41.940 77.320 ;
        RECT 43.030 77.275 43.320 77.320 ;
      LAYER met1 ;
        RECT 56.790 77.460 57.110 77.520 ;
        RECT 59.090 77.460 59.410 77.520 ;
        RECT 73.440 77.460 73.580 77.615 ;
        RECT 56.790 77.320 73.580 77.460 ;
      LAYER met1 ;
        RECT 73.830 77.460 74.120 77.505 ;
        RECT 76.150 77.460 76.440 77.505 ;
        RECT 77.530 77.460 77.820 77.505 ;
        RECT 73.830 77.320 77.820 77.460 ;
      LAYER met1 ;
        RECT 56.790 77.260 57.110 77.320 ;
        RECT 59.090 77.260 59.410 77.320 ;
      LAYER met1 ;
        RECT 73.830 77.275 74.120 77.320 ;
        RECT 76.150 77.275 76.440 77.320 ;
        RECT 77.530 77.275 77.820 77.320 ;
      LAYER met1 ;
        RECT 40.690 67.940 41.010 68.000 ;
        RECT 56.790 67.940 57.110 68.000 ;
        RECT 40.690 67.800 57.110 67.940 ;
        RECT 40.690 67.740 41.010 67.800 ;
        RECT 56.790 67.740 57.110 67.800 ;
        RECT 57.725 67.260 58.015 67.305 ;
        RECT 62.770 67.260 63.090 67.320 ;
        RECT 57.725 67.120 63.090 67.260 ;
        RECT 57.725 67.075 58.015 67.120 ;
        RECT 62.770 67.060 63.090 67.120 ;
      LAYER met1 ;
        RECT 60.950 64.880 61.240 64.925 ;
        RECT 63.270 64.880 63.560 64.925 ;
        RECT 64.650 64.880 64.940 64.925 ;
        RECT 60.950 64.740 64.940 64.880 ;
        RECT 60.950 64.695 61.240 64.740 ;
        RECT 63.270 64.695 63.560 64.740 ;
        RECT 64.650 64.695 64.940 64.740 ;
      LAYER met1 ;
        RECT 60.485 64.200 60.775 64.245 ;
        RECT 60.930 64.200 61.250 64.260 ;
        RECT 61.850 64.200 62.170 64.260 ;
        RECT 60.485 64.060 61.250 64.200 ;
        RECT 61.655 64.060 62.170 64.200 ;
        RECT 60.485 64.015 60.775 64.060 ;
        RECT 60.930 64.000 61.250 64.060 ;
        RECT 61.850 64.000 62.170 64.060 ;
      LAYER met1 ;
        RECT 61.410 63.860 61.700 63.905 ;
        RECT 62.810 63.860 63.100 63.905 ;
        RECT 64.650 63.860 64.940 63.905 ;
        RECT 61.410 63.720 64.940 63.860 ;
        RECT 61.410 63.675 61.700 63.720 ;
        RECT 62.810 63.675 63.100 63.720 ;
        RECT 64.650 63.675 64.940 63.720 ;
        RECT 41.630 62.160 41.920 62.205 ;
        RECT 43.030 62.160 43.320 62.205 ;
        RECT 44.870 62.160 45.160 62.205 ;
        RECT 41.630 62.020 45.160 62.160 ;
        RECT 41.630 61.975 41.920 62.020 ;
        RECT 43.030 61.975 43.320 62.020 ;
        RECT 44.870 61.975 45.160 62.020 ;
        RECT 69.690 62.160 69.980 62.205 ;
        RECT 71.090 62.160 71.380 62.205 ;
        RECT 72.930 62.160 73.220 62.205 ;
        RECT 69.690 62.020 73.220 62.160 ;
        RECT 69.690 61.975 69.980 62.020 ;
        RECT 71.090 61.975 71.380 62.020 ;
        RECT 72.930 61.975 73.220 62.020 ;
      LAYER met1 ;
        RECT 40.690 61.820 41.010 61.880 ;
        RECT 60.010 61.820 60.330 61.880 ;
        RECT 40.495 61.680 41.010 61.820 ;
        RECT 59.815 61.680 60.330 61.820 ;
        RECT 40.690 61.620 41.010 61.680 ;
        RECT 60.010 61.620 60.330 61.680 ;
        RECT 42.070 61.480 42.390 61.540 ;
        RECT 41.875 61.340 42.390 61.480 ;
        RECT 42.070 61.280 42.390 61.340 ;
        RECT 56.790 61.480 57.110 61.540 ;
        RECT 68.765 61.480 69.055 61.525 ;
        RECT 70.130 61.480 70.450 61.540 ;
        RECT 56.790 61.340 69.055 61.480 ;
        RECT 69.935 61.340 70.450 61.480 ;
        RECT 56.790 61.280 57.110 61.340 ;
        RECT 68.765 61.295 69.055 61.340 ;
        RECT 70.130 61.280 70.450 61.340 ;
      LAYER met1 ;
        RECT 41.170 61.140 41.460 61.185 ;
        RECT 43.490 61.140 43.780 61.185 ;
        RECT 44.870 61.140 45.160 61.185 ;
        RECT 41.170 61.000 45.160 61.140 ;
        RECT 41.170 60.955 41.460 61.000 ;
        RECT 43.490 60.955 43.780 61.000 ;
        RECT 44.870 60.955 45.160 61.000 ;
        RECT 69.230 61.140 69.520 61.185 ;
        RECT 71.550 61.140 71.840 61.185 ;
        RECT 72.930 61.140 73.220 61.185 ;
        RECT 69.230 61.000 73.220 61.140 ;
        RECT 69.230 60.955 69.520 61.000 ;
        RECT 71.550 60.955 71.840 61.000 ;
        RECT 72.930 60.955 73.220 61.000 ;
      LAYER met1 ;
        RECT 60.945 60.800 61.235 60.845 ;
        RECT 63.690 60.800 64.010 60.860 ;
        RECT 60.945 60.660 64.010 60.800 ;
        RECT 60.945 60.615 61.235 60.660 ;
        RECT 63.690 60.600 64.010 60.660 ;
        RECT 37.930 59.780 38.250 59.840 ;
        RECT 61.850 59.780 62.170 59.840 ;
        RECT 65.085 59.780 65.375 59.825 ;
        RECT 37.930 59.640 38.620 59.780 ;
        RECT 37.930 59.580 38.250 59.640 ;
        RECT 38.480 59.440 38.620 59.640 ;
        RECT 61.850 59.640 65.375 59.780 ;
        RECT 61.850 59.580 62.170 59.640 ;
        RECT 65.085 59.595 65.375 59.640 ;
        RECT 60.010 59.440 60.330 59.500 ;
        RECT 38.480 59.300 60.330 59.440 ;
        RECT 38.480 58.805 38.620 59.300 ;
        RECT 60.010 59.240 60.330 59.300 ;
        RECT 40.705 59.100 40.995 59.145 ;
        RECT 42.070 59.100 42.390 59.160 ;
        RECT 40.705 58.960 42.390 59.100 ;
        RECT 40.705 58.915 40.995 58.960 ;
        RECT 42.070 58.900 42.390 58.960 ;
        RECT 38.405 58.575 38.695 58.805 ;
        RECT 63.690 58.760 64.010 58.820 ;
        RECT 63.495 58.620 64.010 58.760 ;
        RECT 63.690 58.560 64.010 58.620 ;
        RECT 67.845 56.720 68.135 56.765 ;
        RECT 70.130 56.720 70.450 56.780 ;
        RECT 67.845 56.580 70.450 56.720 ;
        RECT 67.845 56.535 68.135 56.580 ;
        RECT 70.130 56.520 70.450 56.580 ;
        RECT 61.850 56.040 62.170 56.100 ;
        RECT 63.690 56.040 64.010 56.100 ;
        RECT 65.085 56.040 65.375 56.085 ;
        RECT 61.850 55.900 65.375 56.040 ;
        RECT 61.850 55.840 62.170 55.900 ;
        RECT 63.690 55.840 64.010 55.900 ;
        RECT 65.085 55.855 65.375 55.900 ;
        RECT 62.770 54.000 63.090 54.060 ;
        RECT 62.575 53.860 63.090 54.000 ;
        RECT 62.770 53.800 63.090 53.860 ;
      LAYER met1 ;
        RECT 61.870 51.280 62.160 51.325 ;
        RECT 63.270 51.280 63.560 51.325 ;
        RECT 65.110 51.280 65.400 51.325 ;
        RECT 61.870 51.140 65.400 51.280 ;
        RECT 61.870 51.095 62.160 51.140 ;
        RECT 63.270 51.095 63.560 51.140 ;
        RECT 65.110 51.095 65.400 51.140 ;
      LAYER met1 ;
        RECT 60.930 50.940 61.250 51.000 ;
        RECT 60.735 50.800 61.250 50.940 ;
        RECT 60.930 50.740 61.250 50.800 ;
        RECT 62.310 50.600 62.630 50.660 ;
        RECT 62.115 50.460 62.630 50.600 ;
        RECT 62.310 50.400 62.630 50.460 ;
      LAYER met1 ;
        RECT 61.410 50.260 61.700 50.305 ;
        RECT 63.730 50.260 64.020 50.305 ;
        RECT 65.110 50.260 65.400 50.305 ;
        RECT 61.410 50.120 65.400 50.260 ;
        RECT 61.410 50.075 61.700 50.120 ;
        RECT 63.730 50.075 64.020 50.120 ;
        RECT 65.110 50.075 65.400 50.120 ;
      LAYER met1 ;
        RECT 59.565 48.900 59.855 48.945 ;
        RECT 60.930 48.900 61.250 48.960 ;
        RECT 59.565 48.760 61.250 48.900 ;
        RECT 59.565 48.715 59.855 48.760 ;
        RECT 60.930 48.700 61.250 48.760 ;
        RECT 60.485 47.880 60.775 47.925 ;
        RECT 62.770 47.880 63.090 47.940 ;
        RECT 60.485 47.740 63.090 47.880 ;
        RECT 60.485 47.695 60.775 47.740 ;
        RECT 62.770 47.680 63.090 47.740 ;
        RECT 62.310 45.840 62.630 45.900 ;
        RECT 62.115 45.700 62.630 45.840 ;
        RECT 62.310 45.640 62.630 45.700 ;
        RECT 59.550 45.160 59.870 45.220 ;
        RECT 59.355 45.020 59.870 45.160 ;
        RECT 59.550 44.960 59.870 45.020 ;
        RECT 61.850 23.740 62.170 23.800 ;
        RECT 72.905 23.740 73.195 23.785 ;
        RECT 61.850 23.600 73.195 23.740 ;
        RECT 61.850 23.540 62.170 23.600 ;
        RECT 72.905 23.555 73.195 23.600 ;
        RECT 74.285 22.720 74.575 22.765 ;
        RECT 74.730 22.720 75.050 22.780 ;
        RECT 74.285 22.580 75.050 22.720 ;
        RECT 74.285 22.535 74.575 22.580 ;
        RECT 74.730 22.520 75.050 22.580 ;
      LAYER met1 ;
        RECT 54.510 21.360 54.800 21.405 ;
        RECT 56.830 21.360 57.120 21.405 ;
        RECT 58.210 21.360 58.500 21.405 ;
        RECT 54.510 21.220 58.500 21.360 ;
        RECT 54.510 21.175 54.800 21.220 ;
        RECT 56.830 21.175 57.120 21.220 ;
        RECT 58.210 21.175 58.500 21.220 ;
        RECT 73.830 21.360 74.120 21.405 ;
        RECT 76.150 21.360 76.440 21.405 ;
        RECT 77.530 21.360 77.820 21.405 ;
        RECT 73.830 21.220 77.820 21.360 ;
        RECT 73.830 21.175 74.120 21.220 ;
        RECT 76.150 21.175 76.440 21.220 ;
        RECT 77.530 21.175 77.820 21.220 ;
      LAYER met1 ;
        RECT 54.045 21.020 54.335 21.065 ;
        RECT 60.930 21.020 61.250 21.080 ;
        RECT 73.365 21.020 73.655 21.065 ;
        RECT 74.730 21.020 75.050 21.080 ;
        RECT 54.045 20.880 73.655 21.020 ;
        RECT 74.535 20.880 75.050 21.020 ;
        RECT 54.045 20.835 54.335 20.880 ;
        RECT 60.930 20.820 61.250 20.880 ;
        RECT 73.365 20.835 73.655 20.880 ;
        RECT 74.730 20.820 75.050 20.880 ;
        RECT 55.425 20.680 55.715 20.725 ;
        RECT 61.390 20.680 61.710 20.740 ;
        RECT 55.425 20.540 61.710 20.680 ;
        RECT 55.425 20.495 55.715 20.540 ;
        RECT 61.390 20.480 61.710 20.540 ;
      LAYER met1 ;
        RECT 54.970 20.340 55.260 20.385 ;
        RECT 56.370 20.340 56.660 20.385 ;
        RECT 58.210 20.340 58.500 20.385 ;
        RECT 54.970 20.200 58.500 20.340 ;
        RECT 54.970 20.155 55.260 20.200 ;
        RECT 56.370 20.155 56.660 20.200 ;
        RECT 58.210 20.155 58.500 20.200 ;
        RECT 74.290 20.340 74.580 20.385 ;
        RECT 75.690 20.340 75.980 20.385 ;
        RECT 77.530 20.340 77.820 20.385 ;
        RECT 74.290 20.200 77.820 20.340 ;
        RECT 74.290 20.155 74.580 20.200 ;
        RECT 75.690 20.155 75.980 20.200 ;
        RECT 77.530 20.155 77.820 20.200 ;
      LAYER met1 ;
        RECT 59.550 18.300 59.870 18.360 ;
        RECT 60.025 18.300 60.315 18.345 ;
        RECT 59.550 18.160 60.315 18.300 ;
        RECT 59.550 18.100 59.870 18.160 ;
        RECT 60.025 18.115 60.315 18.160 ;
        RECT 61.390 17.280 61.710 17.340 ;
        RECT 61.195 17.140 61.710 17.280 ;
        RECT 61.390 17.080 61.710 17.140 ;
      LAYER via ;
        RECT 64.180 91.200 64.440 91.460 ;
        RECT 63.720 90.860 63.980 91.120 ;
        RECT 59.580 88.820 59.840 89.080 ;
        RECT 63.720 88.820 63.980 89.080 ;
        RECT 37.960 82.360 38.220 82.620 ;
        RECT 37.960 80.320 38.220 80.580 ;
        RECT 40.260 79.980 40.520 80.240 ;
        RECT 40.260 77.940 40.520 78.200 ;
        RECT 63.720 77.940 63.980 78.200 ;
        RECT 40.720 77.600 40.980 77.860 ;
        RECT 56.820 77.260 57.080 77.520 ;
        RECT 59.120 77.260 59.380 77.520 ;
        RECT 40.720 67.740 40.980 68.000 ;
        RECT 56.820 67.740 57.080 68.000 ;
        RECT 62.800 67.060 63.060 67.320 ;
        RECT 60.960 64.000 61.220 64.260 ;
        RECT 61.880 64.000 62.140 64.260 ;
        RECT 40.720 61.620 40.980 61.880 ;
        RECT 60.040 61.620 60.300 61.880 ;
        RECT 42.100 61.280 42.360 61.540 ;
        RECT 56.820 61.280 57.080 61.540 ;
        RECT 70.160 61.280 70.420 61.540 ;
        RECT 63.720 60.600 63.980 60.860 ;
        RECT 37.960 59.580 38.220 59.840 ;
        RECT 61.880 59.580 62.140 59.840 ;
        RECT 60.040 59.240 60.300 59.500 ;
        RECT 42.100 58.900 42.360 59.160 ;
        RECT 63.720 58.560 63.980 58.820 ;
        RECT 70.160 56.520 70.420 56.780 ;
        RECT 61.880 55.840 62.140 56.100 ;
        RECT 63.720 55.840 63.980 56.100 ;
        RECT 62.800 53.800 63.060 54.060 ;
        RECT 60.960 50.740 61.220 51.000 ;
        RECT 62.340 50.400 62.600 50.660 ;
        RECT 60.960 48.700 61.220 48.960 ;
        RECT 62.800 47.680 63.060 47.940 ;
        RECT 62.340 45.640 62.600 45.900 ;
        RECT 59.580 44.960 59.840 45.220 ;
        RECT 61.880 23.540 62.140 23.800 ;
        RECT 74.760 22.520 75.020 22.780 ;
        RECT 60.960 20.820 61.220 21.080 ;
        RECT 74.760 20.820 75.020 21.080 ;
        RECT 61.420 20.480 61.680 20.740 ;
        RECT 59.580 18.100 59.840 18.360 ;
        RECT 61.420 17.080 61.680 17.340 ;
      LAYER met2 ;
        RECT 64.180 91.170 64.440 91.490 ;
        RECT 63.720 90.830 63.980 91.150 ;
        RECT 63.780 89.110 63.920 90.830 ;
        RECT 59.580 88.790 59.840 89.110 ;
        RECT 63.720 88.790 63.980 89.110 ;
        RECT 37.960 82.330 38.220 82.650 ;
        RECT 38.020 80.610 38.160 82.330 ;
        RECT 59.640 81.030 59.780 88.790 ;
        RECT 59.180 80.890 59.780 81.030 ;
        RECT 37.960 80.290 38.220 80.610 ;
        RECT 38.020 59.870 38.160 80.290 ;
        RECT 40.260 79.950 40.520 80.270 ;
        RECT 40.320 78.230 40.460 79.950 ;
        RECT 40.260 77.910 40.520 78.230 ;
        RECT 40.720 77.570 40.980 77.890 ;
        RECT 40.780 68.030 40.920 77.570 ;
        RECT 59.180 77.550 59.320 80.890 ;
        RECT 64.240 78.310 64.380 91.170 ;
        RECT 63.780 78.230 64.380 78.310 ;
        RECT 63.720 78.170 64.380 78.230 ;
        RECT 63.720 77.910 63.980 78.170 ;
        RECT 56.820 77.230 57.080 77.550 ;
        RECT 59.120 77.230 59.380 77.550 ;
        RECT 56.880 68.030 57.020 77.230 ;
        RECT 40.720 67.710 40.980 68.030 ;
        RECT 56.820 67.710 57.080 68.030 ;
        RECT 40.780 61.910 40.920 67.710 ;
        RECT 40.720 61.590 40.980 61.910 ;
        RECT 56.880 61.570 57.020 67.710 ;
        RECT 62.800 67.030 63.060 67.350 ;
        RECT 60.960 63.970 61.220 64.290 ;
        RECT 61.880 63.970 62.140 64.290 ;
        RECT 60.040 61.590 60.300 61.910 ;
        RECT 42.100 61.250 42.360 61.570 ;
        RECT 56.820 61.250 57.080 61.570 ;
        RECT 37.960 59.550 38.220 59.870 ;
        RECT 42.160 59.190 42.300 61.250 ;
        RECT 60.100 59.530 60.240 61.590 ;
        RECT 60.040 59.210 60.300 59.530 ;
        RECT 42.100 58.870 42.360 59.190 ;
        RECT 60.100 51.790 60.240 59.210 ;
        RECT 59.640 51.650 60.240 51.790 ;
        RECT 59.640 45.250 59.780 51.650 ;
        RECT 61.020 51.030 61.160 63.970 ;
        RECT 61.940 59.870 62.080 63.970 ;
        RECT 61.880 59.550 62.140 59.870 ;
        RECT 61.880 55.810 62.140 56.130 ;
        RECT 60.960 50.710 61.220 51.030 ;
        RECT 61.020 48.990 61.160 50.710 ;
        RECT 60.960 48.670 61.220 48.990 ;
        RECT 59.580 44.930 59.840 45.250 ;
        RECT 59.640 18.390 59.780 44.930 ;
        RECT 61.020 21.110 61.160 48.670 ;
        RECT 61.940 23.830 62.080 55.810 ;
        RECT 62.860 54.090 63.000 67.030 ;
        RECT 63.780 60.890 63.920 77.910 ;
        RECT 70.160 61.250 70.420 61.570 ;
        RECT 63.720 60.570 63.980 60.890 ;
        RECT 63.780 58.850 63.920 60.570 ;
        RECT 63.720 58.530 63.980 58.850 ;
        RECT 63.780 56.130 63.920 58.530 ;
        RECT 70.220 56.810 70.360 61.250 ;
        RECT 70.160 56.490 70.420 56.810 ;
        RECT 63.720 55.810 63.980 56.130 ;
        RECT 62.800 53.770 63.060 54.090 ;
        RECT 62.340 50.370 62.600 50.690 ;
        RECT 62.400 45.930 62.540 50.370 ;
        RECT 62.860 47.970 63.000 53.770 ;
        RECT 62.800 47.650 63.060 47.970 ;
        RECT 62.340 45.610 62.600 45.930 ;
        RECT 61.880 23.510 62.140 23.830 ;
        RECT 74.760 22.490 75.020 22.810 ;
        RECT 74.820 21.110 74.960 22.490 ;
        RECT 60.960 20.790 61.220 21.110 ;
        RECT 74.760 20.790 75.020 21.110 ;
        RECT 61.420 20.450 61.680 20.770 ;
        RECT 59.580 18.070 59.840 18.390 ;
        RECT 61.480 17.370 61.620 20.450 ;
        RECT 61.420 17.050 61.680 17.370 ;
  END
END testdesign
END LIBRARY

